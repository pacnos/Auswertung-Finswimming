<?xml version="1.0" encoding="UTF-8"?>
<LENEX version="3.0">
  <CONSTRUCTOR name="EasyWk" version="5.23" registration="">
    <CONTACT name="Bjoern Stickan" internet="http://www.easywk.de" email="info@easywk.de" />
  </CONSTRUCTOR>
  <MEETS>
    <MEET city="Halle (Saale)" course="LCM" name="Sommer Sprint Cup 2023" nation="GER" organizer="Tauchsport / Flossenschwimmen" hostclub="Schwimm und Sportclub Halle" deadline="2023-06-08" timing="AUTOMATIC">
      <CONTACT email="joehoffmann@gmx.de" name="Hoffmann, Jörg" />
      <AGEDATE type="YEAR" value="2023-01-01" />
      <SESSIONS>
        <SESSION number="1" date="2023-06-17" daytime="10:00" officialmeeting="09:30" warmupfrom="08:45">
          <EVENTS>
            <EVENT eventid="1" number="1" gender="X" round="TIM">
              <SWIMSTYLE stroke="APNEA" relaycount="1" distance="50" />
              <FEE value="500" currency="EUR" />
              <HEATS>
                <HEAT heatid="1001" number="1" />
                <HEAT heatid="1002" number="2" />
                <HEAT heatid="1003" number="3" />
                <HEAT heatid="1004" number="4" />
                <HEAT heatid="1005" number="5" />
                <HEAT heatid="1006" number="6" />
                <HEAT heatid="1007" number="7" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="4" agemax="15" agemin="14" name="Kategorie B weiblich">
                  <RANKINGS>
                    <RANKING place="5" resultid="193" />
                    <RANKING place="8" resultid="333" />
                    <RANKING place="4" resultid="495" />
                    <RANKING place="2" resultid="500" />
                    <RANKING place="6" resultid="545" />
                    <RANKING place="3" resultid="570" />
                    <RANKING place="7" resultid="618" />
                    <RANKING place="1" resultid="630" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="17" agemin="16" name="Kategorie A weiblich">
                  <RANKINGS>
                    <RANKING place="5" resultid="86" />
                    <RANKING place="8" resultid="103" />
                    <RANKING place="1" resultid="136" />
                    <RANKING place="2" resultid="296" />
                    <RANKING place="3" resultid="403" />
                    <RANKING place="7" resultid="441" />
                    <RANKING place="6" resultid="527" />
                    <RANKING place="4" resultid="651" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6" agemax="21" agemin="18" name="Junioren weiblich">
                  <RANKINGS>
                    <RANKING place="7" resultid="1" />
                    <RANKING place="5" resultid="13" />
                    <RANKING place="4" resultid="41" />
                    <RANKING place="6" resultid="48" />
                    <RANKING place="3" resultid="59" />
                    <RANKING place="8" resultid="77" />
                    <RANKING place="1" resultid="189" />
                    <RANKING place="2" resultid="381" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7" agemax="25" agemin="22" name="Pre-Master weiblich" />
                <AGEGROUP agegroupid="8" agemax="-1" agemin="26" name="Master weiblich">
                  <RANKINGS>
                    <RANKING place="1" resultid="6" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="12" agemax="15" agemin="14" name="Kategorie B männlich">
                  <RANKINGS>
                    <RANKING place="4" resultid="37" />
                    <RANKING place="2" resultid="228" />
                    <RANKING place="3" resultid="318" />
                    <RANKING place="6" resultid="347" />
                    <RANKING place="1" resultid="470" />
                    <RANKING place="5" resultid="589" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="13" agemax="17" agemin="16" name="Kategorie A männlich">
                  <RANKINGS>
                    <RANKING place="3" resultid="267" />
                    <RANKING place="2" resultid="377" />
                    <RANKING place="1" resultid="420" />
                    <RANKING place="4" resultid="551" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="14" agemax="21" agemin="18" name="Junioren männlich">
                  <RANKINGS>
                    <RANKING place="5" resultid="55" />
                    <RANKING place="4" resultid="322" />
                    <RANKING place="1" resultid="429" />
                    <RANKING place="3" resultid="483" />
                    <RANKING place="2" resultid="514" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15" agemax="25" agemin="22" name="Pre-Master männlich">
                  <RANKINGS>
                    <RANKING place="2" resultid="307" />
                    <RANKING place="1" resultid="537" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="16" agemax="-1" agemin="26" name="Master männlich">
                  <RANKINGS>
                    <RANKING place="2" resultid="26" />
                    <RANKING place="1" resultid="120" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="17" agemax="15" agemin="14" name="Kategorie B weiblich - LM">
                  <RANKINGS>
                    <RANKING place="2" resultid="495" />
                    <RANKING place="1" resultid="500" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="18" agemax="17" agemin="16" name="Kategorie A weiblich - LM">
                  <RANKINGS>
                    <RANKING place="1" resultid="296" />
                    <RANKING place="4" resultid="441" />
                    <RANKING place="3" resultid="527" />
                    <RANKING place="2" resultid="651" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="19" agemax="21" agemin="18" name="Junioren weiblich - LM" />
                <AGEGROUP agegroupid="20" agemax="25" agemin="22" name="Pre-Master weiblich - LM" />
                <AGEGROUP agegroupid="21" agemax="-1" agemin="26" name="Master weiblich - LM" />
                <AGEGROUP agegroupid="22" agemax="15" agemin="14" name="Kategorie B männlich - LM">
                  <RANKINGS>
                    <RANKING place="2" resultid="318" />
                    <RANKING place="1" resultid="470" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="23" agemax="17" agemin="16" name="Kategorie A männlich - LM">
                  <RANKINGS>
                    <RANKING place="1" resultid="267" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="24" agemax="21" agemin="18" name="Junioren männlich - LM">
                  <RANKINGS>
                    <RANKING place="3" resultid="322" />
                    <RANKING place="2" resultid="483" />
                    <RANKING place="1" resultid="514" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="25" agemax="25" agemin="22" name="Pre-Master männlich - LM">
                  <RANKINGS>
                    <RANKING place="1" resultid="307" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="26" agemax="-1" agemin="26" name="Master männlich - LM" />
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="2" number="101" gender="X" round="TIM">
              <SWIMSTYLE stroke="FREE" technique="KICK" relaycount="1" distance="50" />
              <FEE value="500" currency="EUR" />
              <HEATS>
                <HEAT heatid="2001" number="1" />
                <HEAT heatid="2002" number="2" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="8" agemin="0" name="Jg. 2015 u. jünger weiblich">
                  <RANKINGS>
                    <RANKING place="4" resultid="123" />
                    <RANKING place="1" resultid="144" />
                    <RANKING place="3" resultid="373" />
                    <RANKING place="2" resultid="523" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2" agemax="8" agemin="0" name="Jg. 2015 u. jünger männlich">
                  <RANKINGS>
                    <RANKING place="3" resultid="157" />
                    <RANKING place="1" resultid="221" />
                    <RANKING place="2" resultid="243" />
                    <RANKING place="5" resultid="271" />
                    <RANKING place="9" resultid="286" />
                    <RANKING place="8" resultid="303" />
                    <RANKING place="7" resultid="313" />
                    <RANKING place="6" resultid="556" />
                    <RANKING place="4" resultid="601" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3" agemax="8" agemin="0" name="Jg. 2015 u. jünger weiblich - LM">
                  <RANKINGS>
                    <RANKING place="1" resultid="523" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="8" agemin="0" name="Jg. 2015 u. jünger männlich - LM">
                  <RANKINGS>
                    <RANKING place="1" resultid="271" />
                    <RANKING place="4" resultid="286" />
                    <RANKING place="3" resultid="303" />
                    <RANKING place="2" resultid="313" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="3" number="2" gender="X" round="TIM">
              <SWIMSTYLE stroke="SURFACE" relaycount="1" distance="400" />
              <FEE value="500" currency="EUR" />
              <HEATS>
                <HEAT heatid="3001" number="1" />
                <HEAT heatid="3002" number="2" />
                <HEAT heatid="3003" number="3" />
                <HEAT heatid="3004" number="4" />
                <HEAT heatid="3005" number="5" />
                <HEAT heatid="3006" number="6" />
                <HEAT heatid="3007" number="7" />
                <HEAT heatid="3008" number="8" />
                <HEAT heatid="3009" number="9" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="9" agemin="9" name="Kategorie E weiblich">
                  <RANKINGS>
                    <RANKING place="1" resultid="386" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2" agemax="11" agemin="10" name="Kategorie D weiblich">
                  <RANKINGS>
                    <RANKING place="2" resultid="81" />
                    <RANKING place="1" resultid="152" />
                    <RANKING place="4" resultid="160" />
                    <RANKING place="6" resultid="168" />
                    <RANKING place="9" resultid="179" />
                    <RANKING place="5" resultid="184" />
                    <RANKING place="7" resultid="393" />
                    <RANKING place="3" resultid="414" />
                    <RANKING place="8" resultid="487" />
                    <RANKING place="10" resultid="510" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3" agemax="13" agemin="12" name="Kategorie C weiblich">
                  <RANKINGS>
                    <RANKING place="1" resultid="22" />
                    <RANKING place="8" resultid="66" />
                    <RANKING place="3" resultid="70" />
                    <RANKING place="6" resultid="173" />
                    <RANKING place="9" resultid="200" />
                    <RANKING place="7" resultid="232" />
                    <RANKING place="12" resultid="236" />
                    <RANKING place="4" resultid="338" />
                    <RANKING place="5" resultid="351" />
                    <RANKING place="10" resultid="479" />
                    <RANKING place="2" resultid="562" />
                    <RANKING place="11" resultid="574" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="15" agemin="14" name="Kategorie B weiblich">
                  <RANKINGS>
                    <RANKING place="5" resultid="33" />
                    <RANKING place="3" resultid="496" />
                    <RANKING place="2" resultid="501" />
                    <RANKING place="6" resultid="546" />
                    <RANKING place="1" resultid="566" />
                    <RANKING place="7" resultid="586" />
                    <RANKING place="4" resultid="619" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="17" agemin="16" name="Kategorie A weiblich">
                  <RANKINGS>
                    <RANKING place="3" resultid="406" />
                    <RANKING place="1" resultid="424" />
                    <RANKING place="2" resultid="442" />
                    <RANKING place="4" resultid="578" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6" agemax="21" agemin="18" name="Junioren weiblich">
                  <RANKINGS>
                    <RANKING place="1" resultid="2" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7" agemax="25" agemin="22" name="Pre-Master weiblich" />
                <AGEGROUP agegroupid="8" agemax="-1" agemin="26" name="Master weiblich">
                  <RANKINGS>
                    <RANKING place="1" resultid="7" />
                    <RANKING place="3" resultid="109" />
                    <RANKING place="2" resultid="427" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9" agemax="9" agemin="9" name="Kategorie E männlich">
                  <RANKINGS>
                    <RANKING place="2" resultid="245" />
                    <RANKING place="1" resultid="437" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10" agemax="11" agemin="10" name="Kategorie D männlich">
                  <RANKINGS>
                    <RANKING place="2" resultid="250" />
                    <RANKING place="4" resultid="446" />
                    <RANKING place="3" resultid="454" />
                    <RANKING place="1" resultid="519" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11" agemax="13" agemin="12" name="Kategorie C männlich">
                  <RANKINGS>
                    <RANKING place="6" resultid="126" />
                    <RANKING place="5" resultid="163" />
                    <RANKING place="4" resultid="282" />
                    <RANKING place="1" resultid="355" />
                    <RANKING place="2" resultid="433" />
                    <RANKING place="3" resultid="614" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="12" agemax="15" agemin="14" name="Kategorie B männlich">
                  <RANKINGS>
                    <RANKING place="6" resultid="204" />
                    <RANKING place="3" resultid="229" />
                    <RANKING place="2" resultid="275" />
                    <RANKING place="7" resultid="348" />
                    <RANKING place="1" resultid="471" />
                    <RANKING place="4" resultid="506" />
                    <RANKING place="8" resultid="532" />
                    <RANKING place="5" resultid="590" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="13" agemax="17" agemin="16" name="Kategorie A männlich">
                  <RANKINGS>
                    <RANKING place="1" resultid="552" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="14" agemax="21" agemin="18" name="Junioren männlich" />
                <AGEGROUP agegroupid="15" agemax="25" agemin="22" name="Pre-Master männlich" />
                <AGEGROUP agegroupid="16" agemax="-1" agemin="26" name="Master männlich" />
                <AGEGROUP agegroupid="17" agemax="9" agemin="9" name="Kategorie E weiblich - LM" />
                <AGEGROUP agegroupid="18" agemax="11" agemin="10" name="Kategorie D weiblich - LM">
                  <RANKINGS>
                    <RANKING place="1" resultid="487" />
                    <RANKING place="2" resultid="510" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="19" agemax="13" agemin="12" name="Kategorie C weiblich - LM">
                  <RANKINGS>
                    <RANKING place="1" resultid="479" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="20" agemax="15" agemin="14" name="Kategorie B weiblich - LM">
                  <RANKINGS>
                    <RANKING place="2" resultid="496" />
                    <RANKING place="1" resultid="501" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="21" agemax="17" agemin="16" name="Kategorie A weiblich - LM">
                  <RANKINGS>
                    <RANKING place="1" resultid="442" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="22" agemax="21" agemin="18" name="Junioren weiblich - LM" />
                <AGEGROUP agegroupid="23" agemax="25" agemin="22" name="Pre-Master weiblich - LM" />
                <AGEGROUP agegroupid="24" agemax="-1" agemin="26" name="Master weiblich - LM" />
                <AGEGROUP agegroupid="25" agemax="9" agemin="9" name="Kategorie E männlich - LM">
                  <RANKINGS>
                    <RANKING place="1" resultid="437" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="26" agemax="11" agemin="10" name="Kategorie D männlich - LM">
                  <RANKINGS>
                    <RANKING place="3" resultid="446" />
                    <RANKING place="2" resultid="454" />
                    <RANKING place="1" resultid="519" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="27" agemax="13" agemin="12" name="Kategorie C männlich - LM">
                  <RANKINGS>
                    <RANKING place="2" resultid="282" />
                    <RANKING place="1" resultid="433" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="28" agemax="15" agemin="14" name="Kategorie B männlich - LM">
                  <RANKINGS>
                    <RANKING place="2" resultid="275" />
                    <RANKING place="1" resultid="471" />
                    <RANKING place="3" resultid="506" />
                    <RANKING place="4" resultid="532" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="29" agemax="17" agemin="16" name="Kategorie A männlich - LM" />
                <AGEGROUP agegroupid="30" agemax="21" agemin="18" name="Junioren männlich - LM" />
                <AGEGROUP agegroupid="31" agemax="25" agemin="22" name="Pre-Master männlich - LM" />
                <AGEGROUP agegroupid="32" agemax="-1" agemin="26" name="Master männlich - LM" />
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="4" number="102" gender="X" round="TIM">
              <SWIMSTYLE stroke="APNEA" relaycount="1" distance="25" />
              <FEE value="500" currency="EUR" />
              <HEATS>
                <HEAT heatid="4001" number="1" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="8" agemin="0" name="Jg. 2015 u. jünger weiblich">
                  <RANKINGS>
                    <RANKING place="2" resultid="145" />
                    <RANKING place="1" resultid="524" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2" agemax="8" agemin="0" name="Jg. 2015 u. jünger männlich">
                  <RANKINGS>
                    <RANKING place="1" resultid="222" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3" agemax="8" agemin="0" name="Jg. 2015 u. jünger weiblich - LM">
                  <RANKINGS>
                    <RANKING place="1" resultid="524" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="8" agemin="0" name="Jg. 2015 u. jünger männlich - LM" />
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="5" number="3" gender="X" round="PRE">
              <SWIMSTYLE stroke="SURFACE" relaycount="1" distance="100" />
              <FEE value="500" currency="EUR" />
              <HEATS>
                <HEAT heatid="5001" number="1" />
                <HEAT heatid="5002" number="2" />
                <HEAT heatid="5003" number="3" />
                <HEAT heatid="5004" number="4" />
                <HEAT heatid="5005" number="5" />
                <HEAT heatid="5006" number="6" />
                <HEAT heatid="5007" number="7" />
                <HEAT heatid="5008" number="8" />
                <HEAT heatid="5009" number="9" />
                <HEAT heatid="5010" number="10" />
                <HEAT heatid="5011" number="11" />
                <HEAT heatid="5012" number="12" />
                <HEAT heatid="5013" number="13" />
                <HEAT heatid="5014" number="14" />
                <HEAT heatid="5015" number="15" />
                <HEAT heatid="5016" number="16" />
                <HEAT heatid="5017" number="17" />
                <HEAT heatid="5018" number="18" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="9" agemin="9" name="Kategorie E weiblich">
                  <RANKINGS>
                    <RANKING place="3" resultid="148" />
                    <RANKING place="4" resultid="214" />
                    <RANKING place="1" resultid="387" />
                    <RANKING place="2" resultid="458" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2" agemax="11" agemin="10" name="Kategorie D weiblich">
                  <RANKINGS>
                    <RANKING place="4" resultid="82" />
                    <RANKING place="9" resultid="93" />
                    <RANKING place="17" resultid="140" />
                    <RANKING place="2" resultid="153" />
                    <RANKING place="6" resultid="161" />
                    <RANKING place="8" resultid="169" />
                    <RANKING place="7" resultid="180" />
                    <RANKING place="14" resultid="185" />
                    <RANKING place="19" resultid="304" />
                    <RANKING place="18" resultid="394" />
                    <RANKING place="15" resultid="410" />
                    <RANKING place="11" resultid="415" />
                    <RANKING place="13" resultid="467" />
                    <RANKING place="10" resultid="488" />
                    <RANKING place="16" resultid="511" />
                    <RANKING place="3" resultid="622" />
                    <RANKING place="5" resultid="626" />
                    <RANKING place="1" resultid="634" />
                    <RANKING place="12" resultid="647" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3" agemax="13" agemin="12" name="Kategorie C weiblich">
                  <RANKINGS>
                    <RANKING place="3" resultid="23" />
                    <RANKING place="2" resultid="63" />
                    <RANKING place="19" resultid="67" />
                    <RANKING place="5" resultid="71" />
                    <RANKING place="13" resultid="99" />
                    <RANKING place="14" resultid="113" />
                    <RANKING place="10" resultid="115" />
                    <RANKING place="8" resultid="174" />
                    <RANKING place="4" resultid="197" />
                    <RANKING place="17" resultid="201" />
                    <RANKING place="12" resultid="233" />
                    <RANKING place="18" resultid="237" />
                    <RANKING place="21" resultid="264" />
                    <RANKING place="9" resultid="331" />
                    <RANKING place="15" resultid="336" />
                    <RANKING place="6" resultid="339" />
                    <RANKING place="11" resultid="344" />
                    <RANKING place="7" resultid="352" />
                    <RANKING place="16" resultid="451" />
                    <RANKING place="23" resultid="480" />
                    <RANKING place="1" resultid="563" />
                    <RANKING place="20" resultid="575" />
                    <RANKING place="22" resultid="606" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="15" agemin="14" name="Kategorie B weiblich">
                  <RANKINGS>
                    <RANKING place="9" resultid="34" />
                    <RANKING place="5" resultid="194" />
                    <RANKING place="10" resultid="334" />
                    <RANKING place="7" resultid="497" />
                    <RANKING place="2" resultid="502" />
                    <RANKING place="8" resultid="547" />
                    <RANKING place="3" resultid="567" />
                    <RANKING place="4" resultid="572" />
                    <RANKING place="6" resultid="620" />
                    <RANKING place="1" resultid="631" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="17" agemin="16" name="Kategorie A weiblich">
                  <RANKINGS>
                    <RANKING place="4" resultid="87" />
                    <RANKING place="10" resultid="101" />
                    <RANKING place="8" resultid="104" />
                    <RANKING place="9" resultid="118" />
                    <RANKING place="1" resultid="137" />
                    <RANKING place="7" resultid="294" />
                    <RANKING place="2" resultid="297" />
                    <RANKING place="3" resultid="404" />
                    <RANKING place="6" resultid="443" />
                    <RANKING place="5" resultid="529" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6" agemax="21" agemin="18" name="Junioren weiblich">
                  <RANKINGS>
                    <RANKING place="7" resultid="3" />
                    <RANKING place="1" resultid="15" />
                    <RANKING place="5" resultid="49" />
                    <RANKING place="3" resultid="60" />
                    <RANKING place="6" resultid="78" />
                    <RANKING place="2" resultid="190" />
                    <RANKING place="4" resultid="382" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7" agemax="25" agemin="22" name="Pre-Master weiblich">
                  <RANKINGS>
                    <RANKING place="1" resultid="11" />
                    <RANKING place="2" resultid="431" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8" agemax="-1" agemin="26" name="Master weiblich">
                  <RANKINGS>
                    <RANKING place="1" resultid="8" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9" agemax="9" agemin="9" name="Kategorie E männlich">
                  <RANKINGS>
                    <RANKING place="1" resultid="246" />
                    <RANKING place="2" resultid="369" />
                    <RANKING place="4" resultid="438" />
                    <RANKING place="3" resultid="462" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10" agemax="11" agemin="10" name="Kategorie D männlich">
                  <RANKINGS>
                    <RANKING place="1" resultid="251" />
                    <RANKING place="7" resultid="261" />
                    <RANKING place="5" resultid="327" />
                    <RANKING place="4" resultid="447" />
                    <RANKING place="3" resultid="455" />
                    <RANKING place="2" resultid="520" />
                    <RANKING place="6" resultid="541" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11" agemax="13" agemin="12" name="Kategorie C männlich">
                  <RANKINGS>
                    <RANKING place="7" resultid="29" />
                    <RANKING place="9" resultid="107" />
                    <RANKING place="10" resultid="127" />
                    <RANKING place="6" resultid="164" />
                    <RANKING place="4" resultid="283" />
                    <RANKING place="8" resultid="324" />
                    <RANKING place="3" resultid="356" />
                    <RANKING place="11" resultid="391" />
                    <RANKING place="1" resultid="593" />
                    <RANKING place="2" resultid="597" />
                    <RANKING place="5" resultid="615" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="12" agemax="15" agemin="14" name="Kategorie B männlich">
                  <RANKINGS>
                    <RANKING place="4" resultid="38" />
                    <RANKING place="9" resultid="45" />
                    <RANKING place="10" resultid="74" />
                    <RANKING place="11" resultid="95" />
                    <RANKING place="2" resultid="211" />
                    <RANKING place="3" resultid="276" />
                    <RANKING place="5" resultid="319" />
                    <RANKING place="8" resultid="349" />
                    <RANKING place="1" resultid="472" />
                    <RANKING place="6" resultid="507" />
                    <RANKING place="7" resultid="533" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="13" agemax="17" agemin="16" name="Kategorie A männlich">
                  <RANKINGS>
                    <RANKING place="3" resultid="268" />
                    <RANKING place="2" resultid="378" />
                    <RANKING place="1" resultid="421" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="14" agemax="21" agemin="18" name="Junioren männlich">
                  <RANKINGS>
                    <RANKING place="2" resultid="56" />
                    <RANKING place="1" resultid="484" />
                    <RANKING place="3" resultid="492" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15" agemax="25" agemin="22" name="Pre-Master männlich">
                  <RANKINGS>
                    <RANKING place="2" resultid="308" />
                    <RANKING place="3" resultid="315" />
                    <RANKING place="1" resultid="538" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="16" agemax="-1" agemin="26" name="Master männlich">
                  <RANKINGS>
                    <RANKING place="1" resultid="27" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="17" agemax="9" agemin="9" name="Kategorie E weiblich - LM">
                  <RANKINGS>
                    <RANKING place="1" resultid="458" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="18" agemax="11" agemin="10" name="Kategorie D weiblich - LM">
                  <RANKINGS>
                    <RANKING place="4" resultid="304" />
                    <RANKING place="2" resultid="467" />
                    <RANKING place="1" resultid="488" />
                    <RANKING place="3" resultid="511" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="19" agemax="13" agemin="12" name="Kategorie C weiblich - LM">
                  <RANKINGS>
                    <RANKING place="2" resultid="264" />
                    <RANKING place="1" resultid="451" />
                    <RANKING place="3" resultid="480" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="20" agemax="15" agemin="14" name="Kategorie B weiblich - LM">
                  <RANKINGS>
                    <RANKING place="2" resultid="497" />
                    <RANKING place="1" resultid="502" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="21" agemax="17" agemin="16" name="Kategorie A weiblich - LM">
                  <RANKINGS>
                    <RANKING place="4" resultid="294" />
                    <RANKING place="1" resultid="297" />
                    <RANKING place="3" resultid="443" />
                    <RANKING place="2" resultid="529" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="22" agemax="21" agemin="18" name="Junioren weiblich - LM" />
                <AGEGROUP agegroupid="23" agemax="25" agemin="22" name="Pre-Master weiblich - LM" />
                <AGEGROUP agegroupid="24" agemax="-1" agemin="26" name="Master weiblich - LM" />
                <AGEGROUP agegroupid="25" agemax="9" agemin="9" name="Kategorie E männlich - LM">
                  <RANKINGS>
                    <RANKING place="2" resultid="438" />
                    <RANKING place="1" resultid="462" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="26" agemax="11" agemin="10" name="Kategorie D männlich - LM">
                  <RANKINGS>
                    <RANKING place="5" resultid="261" />
                    <RANKING place="4" resultid="327" />
                    <RANKING place="3" resultid="447" />
                    <RANKING place="2" resultid="455" />
                    <RANKING place="1" resultid="520" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="27" agemax="13" agemin="12" name="Kategorie C männlich - LM">
                  <RANKINGS>
                    <RANKING place="1" resultid="283" />
                    <RANKING place="2" resultid="324" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="28" agemax="15" agemin="14" name="Kategorie B männlich - LM">
                  <RANKINGS>
                    <RANKING place="2" resultid="276" />
                    <RANKING place="3" resultid="319" />
                    <RANKING place="1" resultid="472" />
                    <RANKING place="4" resultid="507" />
                    <RANKING place="5" resultid="533" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="29" agemax="17" agemin="16" name="Kategorie A männlich - LM">
                  <RANKINGS>
                    <RANKING place="1" resultid="268" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="30" agemax="21" agemin="18" name="Junioren männlich - LM">
                  <RANKINGS>
                    <RANKING place="1" resultid="484" />
                    <RANKING place="2" resultid="492" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="31" agemax="25" agemin="22" name="Pre-Master männlich - LM">
                  <RANKINGS>
                    <RANKING place="1" resultid="308" />
                    <RANKING place="2" resultid="315" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="32" agemax="-1" agemin="26" name="Master männlich - LM" />
                <AGEGROUP agegroupid="33" agemax="8" agemin="0" name="Jg. 2015 u. jünger">
                  <RANKINGS>
                    <RANKING place="3" resultid="638" />
                    <RANKING place="2" resultid="641" />
                    <RANKING place="1" resultid="643" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="6" number="4" gender="X" round="TIM">
              <SWIMSTYLE stroke="IMMERSION" technique="DIVE" relaycount="1" distance="400" />
              <FEE value="500" currency="EUR" />
              <HEATS>
                <HEAT heatid="6001" number="1" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="9" agemin="9" name="Kategorie E weiblich" />
                <AGEGROUP agegroupid="2" agemax="11" agemin="10" name="Kategorie D weiblich" />
                <AGEGROUP agegroupid="3" agemax="13" agemin="12" name="Kategorie C weiblich" />
                <AGEGROUP agegroupid="4" agemax="15" agemin="14" name="Kategorie B weiblich" />
                <AGEGROUP agegroupid="5" agemax="17" agemin="16" name="Kategorie A weiblich">
                  <RANKINGS>
                    <RANKING place="1" resultid="88" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6" agemax="21" agemin="18" name="Junioren weiblich">
                  <RANKINGS>
                    <RANKING place="1" resultid="43" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7" agemax="25" agemin="22" name="Pre-Master weiblich" />
                <AGEGROUP agegroupid="8" agemax="-1" agemin="26" name="Master weiblich">
                  <RANKINGS>
                    <RANKING place="1" resultid="110" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9" agemax="9" agemin="9" name="Kategorie E männlich" />
                <AGEGROUP agegroupid="10" agemax="11" agemin="10" name="Kategorie D männlich" />
                <AGEGROUP agegroupid="11" agemax="13" agemin="12" name="Kategorie C männlich" />
                <AGEGROUP agegroupid="12" agemax="15" agemin="14" name="Kategorie B männlich">
                  <RANKINGS>
                    <RANKING place="1" resultid="230" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="13" agemax="17" agemin="16" name="Kategorie A männlich">
                  <RANKINGS>
                    <RANKING place="1" resultid="553" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="14" agemax="21" agemin="18" name="Junioren männlich" />
                <AGEGROUP agegroupid="15" agemax="25" agemin="22" name="Pre-Master männlich" />
                <AGEGROUP agegroupid="16" agemax="-1" agemin="26" name="Master männlich" />
                <AGEGROUP agegroupid="17" agemax="9" agemin="9" name="Kategorie E weiblich - LM" />
                <AGEGROUP agegroupid="18" agemax="11" agemin="10" name="Kategorie D weiblich - LM" />
                <AGEGROUP agegroupid="19" agemax="13" agemin="12" name="Kategorie C weiblich - LM" />
                <AGEGROUP agegroupid="20" agemax="15" agemin="14" name="Kategorie B weiblich - LM" />
                <AGEGROUP agegroupid="21" agemax="17" agemin="16" name="Kategorie A weiblich - LM" />
                <AGEGROUP agegroupid="22" agemax="21" agemin="18" name="Junioren weiblich - LM" />
                <AGEGROUP agegroupid="23" agemax="25" agemin="22" name="Pre-Master weiblich - LM" />
                <AGEGROUP agegroupid="24" agemax="-1" agemin="26" name="Master weiblich - LM" />
                <AGEGROUP agegroupid="25" agemax="9" agemin="9" name="Kategorie E männlich - LM" />
                <AGEGROUP agegroupid="26" agemax="11" agemin="10" name="Kategorie D männlich - LM" />
                <AGEGROUP agegroupid="27" agemax="13" agemin="12" name="Kategorie C männlich - LM" />
                <AGEGROUP agegroupid="28" agemax="15" agemin="14" name="Kategorie B männlich - LM" />
                <AGEGROUP agegroupid="29" agemax="17" agemin="16" name="Kategorie A männlich - LM" />
                <AGEGROUP agegroupid="30" agemax="21" agemin="18" name="Junioren männlich - LM" />
                <AGEGROUP agegroupid="31" agemax="25" agemin="22" name="Pre-Master männlich - LM" />
                <AGEGROUP agegroupid="32" agemax="-1" agemin="26" name="Master männlich - LM" />
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="7" number="103" gender="X" round="TIM">
              <SWIMSTYLE stroke="UNKNOWN" relaycount="1" distance="50" />
              <FEE value="500" currency="EUR" />
              <HEATS>
                <HEAT heatid="7001" number="1" />
                <HEAT heatid="7002" number="2" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="8" agemin="0" name="Jg. 2015 u. jünger weiblich">
                  <RANKINGS>
                    <RANKING place="4" resultid="124" />
                    <RANKING place="2" resultid="146" />
                    <RANKING place="3" resultid="375" />
                    <RANKING place="1" resultid="525" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2" agemax="8" agemin="0" name="Jg. 2015 u. jünger männlich">
                  <RANKINGS>
                    <RANKING place="3" resultid="158" />
                    <RANKING place="1" resultid="223" />
                    <RANKING place="2" resultid="244" />
                    <RANKING place="4" resultid="557" />
                    <RANKING place="5" resultid="603" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3" agemax="8" agemin="0" name="Jg. 2015 u. jünger weiblich - LM">
                  <RANKINGS>
                    <RANKING place="1" resultid="525" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="8" agemin="0" name="Jg. 2015 u. jünger männlich - LM" />
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="8" number="5" gender="X" round="TIM">
              <SWIMSTYLE stroke="FLY" technique="KICK" relaycount="1" distance="50" />
              <FEE value="500" currency="EUR" />
              <HEATS>
                <HEAT heatid="8001" number="1" />
                <HEAT heatid="8002" number="2" />
                <HEAT heatid="8003" number="3" />
                <HEAT heatid="8004" number="4" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="9" agemin="9" name="Kategorie E weiblich">
                  <RANKINGS>
                    <RANKING place="5" resultid="52" />
                    <RANKING place="4" resultid="149" />
                    <RANKING place="3" resultid="301" />
                    <RANKING place="1" resultid="388" />
                    <RANKING place="2" resultid="459" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2" agemax="11" agemin="10" name="Kategorie D weiblich">
                  <RANKINGS>
                    <RANKING place="4" resultid="83" />
                    <RANKING place="13" resultid="141" />
                    <RANKING place="2" resultid="154" />
                    <RANKING place="12" resultid="162" />
                    <RANKING place="6" resultid="170" />
                    <RANKING place="5" resultid="181" />
                    <RANKING place="9" resultid="186" />
                    <RANKING place="14" resultid="305" />
                    <RANKING place="11" resultid="395" />
                    <RANKING place="10" resultid="411" />
                    <RANKING place="8" resultid="416" />
                    <RANKING place="3" resultid="623" />
                    <RANKING place="7" resultid="627" />
                    <RANKING place="1" resultid="635" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9" agemax="9" agemin="9" name="Kategorie E männlich">
                  <RANKINGS>
                    <RANKING place="2" resultid="247" />
                    <RANKING place="3" resultid="370" />
                    <RANKING place="1" resultid="463" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10" agemax="11" agemin="10" name="Kategorie D männlich">
                  <RANKINGS>
                    <RANKING place="1" resultid="252" />
                    <RANKING place="5" resultid="262" />
                    <RANKING place="3" resultid="280" />
                    <RANKING place="2" resultid="328" />
                    <RANKING place="4" resultid="542" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11" agemax="9" agemin="9" name="Kategorie E weiblich - LM">
                  <RANKINGS>
                    <RANKING place="2" resultid="301" />
                    <RANKING place="1" resultid="459" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="12" agemax="11" agemin="10" name="Kategorie D weiblich - LM">
                  <RANKINGS>
                    <RANKING place="1" resultid="305" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="13" agemax="9" agemin="9" name="Kategorie E männlich - LM">
                  <RANKINGS>
                    <RANKING place="1" resultid="463" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="14" agemax="11" agemin="10" name="Kategorie D männlich - LM">
                  <RANKINGS>
                    <RANKING place="3" resultid="262" />
                    <RANKING place="2" resultid="280" />
                    <RANKING place="1" resultid="328" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="9" number="6" gender="X" round="FIN">
              <SWIMSTYLE stroke="UNKNOWN" relaycount="3" distance="50" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="9" agemin="9" name="Kategorie E weiblich" />
                <AGEGROUP agegroupid="2" agemax="11" agemin="10" name="Kategorie D weiblich" />
                <AGEGROUP agegroupid="3" agemax="13" agemin="12" name="Kategorie C weiblich" />
                <AGEGROUP agegroupid="4" agemax="15" agemin="14" name="Kategorie B weiblich" />
                <AGEGROUP agegroupid="5" agemax="17" agemin="16" name="Kategorie A weiblich" />
                <AGEGROUP agegroupid="6" agemax="21" agemin="18" name="Junioren weiblich" />
                <AGEGROUP agegroupid="7" agemax="25" agemin="22" name="Pre-Master weiblich" />
                <AGEGROUP agegroupid="8" agemax="-1" agemin="26" name="Master weiblich" />
                <AGEGROUP agegroupid="9" agemax="9" agemin="9" name="Kategorie E männlich" />
                <AGEGROUP agegroupid="10" agemax="11" agemin="10" name="Kategorie D männlich" />
                <AGEGROUP agegroupid="11" agemax="13" agemin="12" name="Kategorie C männlich" />
                <AGEGROUP agegroupid="12" agemax="15" agemin="14" name="Kategorie B männlich" />
                <AGEGROUP agegroupid="13" agemax="17" agemin="16" name="Kategorie A männlich" />
                <AGEGROUP agegroupid="14" agemax="21" agemin="18" name="Junioren männlich" />
                <AGEGROUP agegroupid="15" agemax="25" agemin="22" name="Pre-Master männlich" />
                <AGEGROUP agegroupid="16" agemax="-1" agemin="26" name="Master männlich" />
                <AGEGROUP agegroupid="17" agemax="9" agemin="9" name="Kategorie E weiblich - LM" />
                <AGEGROUP agegroupid="18" agemax="11" agemin="10" name="Kategorie D weiblich - LM" />
                <AGEGROUP agegroupid="19" agemax="13" agemin="12" name="Kategorie C weiblich - LM" />
                <AGEGROUP agegroupid="20" agemax="15" agemin="14" name="Kategorie B weiblich - LM" />
                <AGEGROUP agegroupid="21" agemax="17" agemin="16" name="Kategorie A weiblich - LM" />
                <AGEGROUP agegroupid="22" agemax="21" agemin="18" name="Junioren weiblich - LM" />
                <AGEGROUP agegroupid="23" agemax="25" agemin="22" name="Pre-Master weiblich - LM" />
                <AGEGROUP agegroupid="24" agemax="-1" agemin="26" name="Master weiblich - LM" />
                <AGEGROUP agegroupid="25" agemax="9" agemin="9" name="Kategorie E männlich - LM" />
                <AGEGROUP agegroupid="26" agemax="11" agemin="10" name="Kategorie D männlich - LM" />
                <AGEGROUP agegroupid="27" agemax="13" agemin="12" name="Kategorie C männlich - LM" />
                <AGEGROUP agegroupid="28" agemax="15" agemin="14" name="Kategorie B männlich - LM" />
                <AGEGROUP agegroupid="29" agemax="17" agemin="16" name="Kategorie A männlich - LM" />
                <AGEGROUP agegroupid="30" agemax="21" agemin="18" name="Junioren männlich - LM" />
                <AGEGROUP agegroupid="31" agemax="25" agemin="22" name="Pre-Master männlich - LM" />
                <AGEGROUP agegroupid="32" agemax="-1" agemin="26" name="Master männlich - LM" />
              </AGEGROUPS>
            </EVENT>
          </EVENTS>
        </SESSION>
        <SESSION number="2" date="2023-06-17" daytime="00:45">
          <EVENTS>
            <EVENT eventid="10" number="7" gender="X" round="TIM">
              <SWIMSTYLE stroke="SURFACE" relaycount="1" distance="50" />
              <FEE value="500" currency="EUR" />
              <HEATS>
                <HEAT heatid="10001" number="1" />
                <HEAT heatid="10002" number="2" />
                <HEAT heatid="10003" number="3" />
                <HEAT heatid="10004" number="4" />
                <HEAT heatid="10005" number="5" />
                <HEAT heatid="10006" number="6" />
                <HEAT heatid="10007" number="7" />
                <HEAT heatid="10008" number="8" />
                <HEAT heatid="10009" number="9" />
                <HEAT heatid="10010" number="10" />
                <HEAT heatid="10011" number="11" />
                <HEAT heatid="10012" number="12" />
                <HEAT heatid="10013" number="13" />
                <HEAT heatid="10014" number="14" />
                <HEAT heatid="10015" number="15" />
                <HEAT heatid="10016" number="16" />
                <HEAT heatid="10017" number="17" />
                <HEAT heatid="10018" number="18" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="9" agemin="9" name="Kategorie E weiblich">
                  <RANKINGS>
                    <RANKING place="3" resultid="53" />
                    <RANKING place="5" resultid="150" />
                    <RANKING place="6" resultid="216" />
                    <RANKING place="2" resultid="302" />
                    <RANKING place="1" resultid="389" />
                    <RANKING place="4" resultid="460" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2" agemax="11" agemin="10" name="Kategorie D weiblich">
                  <RANKINGS>
                    <RANKING place="9" resultid="84" />
                    <RANKING place="14" resultid="142" />
                    <RANKING place="2" resultid="155" />
                    <RANKING place="7" resultid="171" />
                    <RANKING place="8" resultid="182" />
                    <RANKING place="12" resultid="187" />
                    <RANKING place="15" resultid="306" />
                    <RANKING place="13" resultid="396" />
                    <RANKING place="11" resultid="412" />
                    <RANKING place="10" resultid="417" />
                    <RANKING place="4" resultid="468" />
                    <RANKING place="6" resultid="489" />
                    <RANKING place="3" resultid="624" />
                    <RANKING place="5" resultid="628" />
                    <RANKING place="1" resultid="636" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3" agemax="13" agemin="12" name="Kategorie C weiblich">
                  <RANKINGS>
                    <RANKING place="1" resultid="24" />
                    <RANKING place="3" resultid="64" />
                    <RANKING place="12" resultid="68" />
                    <RANKING place="4" resultid="72" />
                    <RANKING place="17" resultid="100" />
                    <RANKING place="16" resultid="114" />
                    <RANKING place="18" resultid="116" />
                    <RANKING place="6" resultid="175" />
                    <RANKING place="2" resultid="198" />
                    <RANKING place="19" resultid="202" />
                    <RANKING place="14" resultid="234" />
                    <RANKING place="8" resultid="238" />
                    <RANKING place="7" resultid="332" />
                    <RANKING place="13" resultid="337" />
                    <RANKING place="9" resultid="345" />
                    <RANKING place="5" resultid="353" />
                    <RANKING place="10" resultid="362" />
                    <RANKING place="11" resultid="452" />
                    <RANKING place="15" resultid="481" />
                    <RANKING place="20" resultid="576" />
                    <RANKING place="21" resultid="607" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="15" agemin="14" name="Kategorie B weiblich">
                  <RANKINGS>
                    <RANKING place="9" resultid="35" />
                    <RANKING place="6" resultid="195" />
                    <RANKING place="5" resultid="498" />
                    <RANKING place="1" resultid="503" />
                    <RANKING place="8" resultid="548" />
                    <RANKING place="2" resultid="568" />
                    <RANKING place="3" resultid="573" />
                    <RANKING place="10" resultid="587" />
                    <RANKING place="7" resultid="621" />
                    <RANKING place="4" resultid="632" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="17" agemin="16" name="Kategorie A weiblich">
                  <RANKINGS>
                    <RANKING place="3" resultid="89" />
                    <RANKING place="10" resultid="102" />
                    <RANKING place="9" resultid="105" />
                    <RANKING place="8" resultid="119" />
                    <RANKING place="1" resultid="138" />
                    <RANKING place="6" resultid="295" />
                    <RANKING place="2" resultid="298" />
                    <RANKING place="7" resultid="408" />
                    <RANKING place="4" resultid="444" />
                    <RANKING place="5" resultid="530" />
                    <RANKING place="11" resultid="580" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6" agemax="21" agemin="18" name="Junioren weiblich">
                  <RANKINGS>
                    <RANKING place="4" resultid="14" />
                    <RANKING place="5" resultid="50" />
                    <RANKING place="3" resultid="61" />
                    <RANKING place="6" resultid="79" />
                    <RANKING place="2" resultid="191" />
                    <RANKING place="1" resultid="384" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7" agemax="25" agemin="22" name="Pre-Master weiblich">
                  <RANKINGS>
                    <RANKING place="1" resultid="12" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8" agemax="-1" agemin="26" name="Master weiblich">
                  <RANKINGS>
                    <RANKING place="1" resultid="9" />
                    <RANKING place="3" resultid="111" />
                    <RANKING place="2" resultid="428" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9" agemax="9" agemin="9" name="Kategorie E männlich">
                  <RANKINGS>
                    <RANKING place="2" resultid="248" />
                    <RANKING place="5" resultid="312" />
                    <RANKING place="3" resultid="371" />
                    <RANKING place="1" resultid="439" />
                    <RANKING place="4" resultid="464" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10" agemax="11" agemin="10" name="Kategorie D männlich">
                  <RANKINGS>
                    <RANKING place="2" resultid="253" />
                    <RANKING place="8" resultid="263" />
                    <RANKING place="6" resultid="281" />
                    <RANKING place="5" resultid="329" />
                    <RANKING place="1" resultid="448" />
                    <RANKING place="4" resultid="456" />
                    <RANKING place="3" resultid="521" />
                    <RANKING place="7" resultid="543" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11" agemax="13" agemin="12" name="Kategorie C männlich">
                  <RANKINGS>
                    <RANKING place="6" resultid="30" />
                    <RANKING place="7" resultid="108" />
                    <RANKING place="10" resultid="128" />
                    <RANKING place="9" resultid="165" />
                    <RANKING place="3" resultid="284" />
                    <RANKING place="8" resultid="342" />
                    <RANKING place="4" resultid="358" />
                    <RANKING place="11" resultid="392" />
                    <RANKING place="2" resultid="594" />
                    <RANKING place="1" resultid="598" />
                    <RANKING place="5" resultid="616" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="12" agemax="15" agemin="14" name="Kategorie B männlich">
                  <RANKINGS>
                    <RANKING place="4" resultid="39" />
                    <RANKING place="5" resultid="46" />
                    <RANKING place="11" resultid="75" />
                    <RANKING place="6" resultid="206" />
                    <RANKING place="1" resultid="212" />
                    <RANKING place="2" resultid="277" />
                    <RANKING place="3" resultid="320" />
                    <RANKING place="8" resultid="473" />
                    <RANKING place="6" resultid="508" />
                    <RANKING place="9" resultid="534" />
                    <RANKING place="10" resultid="591" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="13" agemax="17" agemin="16" name="Kategorie A männlich">
                  <RANKINGS>
                    <RANKING place="3" resultid="269" />
                    <RANKING place="2" resultid="379" />
                    <RANKING place="1" resultid="422" />
                    <RANKING place="4" resultid="554" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="14" agemax="21" agemin="18" name="Junioren männlich">
                  <RANKINGS>
                    <RANKING place="3" resultid="57" />
                    <RANKING place="4" resultid="323" />
                    <RANKING place="1" resultid="485" />
                    <RANKING place="2" resultid="516" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15" agemax="25" agemin="22" name="Pre-Master männlich">
                  <RANKINGS>
                    <RANKING place="2" resultid="309" />
                    <RANKING place="3" resultid="316" />
                    <RANKING place="1" resultid="539" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="16" agemax="-1" agemin="26" name="Master männlich">
                  <RANKINGS>
                    <RANKING place="2" resultid="28" />
                    <RANKING place="1" resultid="121" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="17" agemax="9" agemin="9" name="Kategorie E weiblich - LM">
                  <RANKINGS>
                    <RANKING place="1" resultid="302" />
                    <RANKING place="2" resultid="460" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="18" agemax="11" agemin="10" name="Kategorie D weiblich - LM">
                  <RANKINGS>
                    <RANKING place="3" resultid="306" />
                    <RANKING place="1" resultid="468" />
                    <RANKING place="2" resultid="489" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="19" agemax="13" agemin="12" name="Kategorie C weiblich - LM">
                  <RANKINGS>
                    <RANKING place="1" resultid="452" />
                    <RANKING place="2" resultid="481" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="20" agemax="15" agemin="14" name="Kategorie B weiblich - LM">
                  <RANKINGS>
                    <RANKING place="2" resultid="498" />
                    <RANKING place="1" resultid="503" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="21" agemax="17" agemin="16" name="Kategorie A weiblich - LM">
                  <RANKINGS>
                    <RANKING place="4" resultid="295" />
                    <RANKING place="1" resultid="298" />
                    <RANKING place="2" resultid="444" />
                    <RANKING place="3" resultid="530" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="22" agemax="21" agemin="18" name="Junioren weiblich - LM" />
                <AGEGROUP agegroupid="23" agemax="25" agemin="22" name="Pre-Master weiblich - LM" />
                <AGEGROUP agegroupid="24" agemax="-1" agemin="26" name="Master weiblich - LM" />
                <AGEGROUP agegroupid="25" agemax="9" agemin="9" name="Kategorie E männlich - LM">
                  <RANKINGS>
                    <RANKING place="3" resultid="312" />
                    <RANKING place="1" resultid="439" />
                    <RANKING place="2" resultid="464" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="26" agemax="11" agemin="10" name="Kategorie D männlich - LM">
                  <RANKINGS>
                    <RANKING place="6" resultid="263" />
                    <RANKING place="5" resultid="281" />
                    <RANKING place="4" resultid="329" />
                    <RANKING place="1" resultid="448" />
                    <RANKING place="3" resultid="456" />
                    <RANKING place="2" resultid="521" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="27" agemax="13" agemin="12" name="Kategorie C männlich - LM">
                  <RANKINGS>
                    <RANKING place="1" resultid="284" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="28" agemax="15" agemin="14" name="Kategorie B männlich - LM">
                  <RANKINGS>
                    <RANKING place="1" resultid="277" />
                    <RANKING place="2" resultid="320" />
                    <RANKING place="4" resultid="473" />
                    <RANKING place="3" resultid="508" />
                    <RANKING place="5" resultid="534" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="29" agemax="17" agemin="16" name="Kategorie A männlich - LM">
                  <RANKINGS>
                    <RANKING place="1" resultid="269" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="30" agemax="21" agemin="18" name="Junioren männlich - LM">
                  <RANKINGS>
                    <RANKING place="3" resultid="323" />
                    <RANKING place="1" resultid="485" />
                    <RANKING place="2" resultid="516" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="31" agemax="25" agemin="22" name="Pre-Master männlich - LM">
                  <RANKINGS>
                    <RANKING place="1" resultid="309" />
                    <RANKING place="2" resultid="316" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="32" agemax="-1" agemin="26" name="Master männlich - LM" />
                <AGEGROUP agegroupid="33" agemax="8" agemin="0" name="Jg. 2015 u. jünger">
                  <RANKINGS>
                    <RANKING place="1" resultid="256" />
                    <RANKING place="3" resultid="642" />
                    <RANKING place="2" resultid="644" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="11" number="104" gender="X" round="TIM">
              <SWIMSTYLE stroke="SURFACE" relaycount="1" distance="50" />
              <FEE value="500" currency="EUR" />
              <HEATS>
                <HEAT heatid="11001" number="1" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="8" agemin="0" name="Jg. 2015 u. jünger weiblich">
                  <RANKINGS>
                    <RANKING place="4" resultid="125" />
                    <RANKING place="3" resultid="147" />
                    <RANKING place="2" resultid="376" />
                    <RANKING place="1" resultid="526" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2" agemax="8" agemin="0" name="Jg. 2015 u. jünger männlich">
                  <RANKINGS>
                    <RANKING place="3" resultid="159" />
                    <RANKING place="2" resultid="558" />
                    <RANKING place="4" resultid="604" />
                    <RANKING place="1" resultid="650" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3" agemax="8" agemin="0" name="Jg. 2015 u. jünger weiblich - LM">
                  <RANKINGS>
                    <RANKING place="1" resultid="526" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="8" agemin="0" name="Jg. 2015 u. jünger männlich - LM" />
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="12" number="8" gender="X" round="TIM">
              <SWIMSTYLE stroke="IMMERSION" technique="DIVE" relaycount="1" distance="100" />
              <FEE value="500" currency="EUR" />
              <HEATS>
                <HEAT heatid="12001" number="1" />
                <HEAT heatid="12002" number="2" />
                <HEAT heatid="12003" number="3" />
                <HEAT heatid="12004" number="4" />
                <HEAT heatid="12005" number="5" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="9" agemin="9" name="Kategorie E weiblich" />
                <AGEGROUP agegroupid="2" agemax="11" agemin="10" name="Kategorie D weiblich" />
                <AGEGROUP agegroupid="3" agemax="13" agemin="12" name="Kategorie C weiblich">
                  <RANKINGS>
                    <RANKING place="3" resultid="176" />
                    <RANKING place="2" resultid="199" />
                    <RANKING place="7" resultid="239" />
                    <RANKING place="5" resultid="341" />
                    <RANKING place="8" resultid="346" />
                    <RANKING place="4" resultid="354" />
                    <RANKING place="6" resultid="363" />
                    <RANKING place="1" resultid="565" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="15" agemin="14" name="Kategorie B weiblich">
                  <RANKINGS>
                    <RANKING place="2" resultid="196" />
                    <RANKING place="5" resultid="335" />
                    <RANKING place="3" resultid="549" />
                    <RANKING place="4" resultid="588" />
                    <RANKING place="1" resultid="633" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="17" agemin="16" name="Kategorie A weiblich">
                  <RANKINGS>
                    <RANKING place="2" resultid="90" />
                    <RANKING place="4" resultid="106" />
                    <RANKING place="1" resultid="139" />
                    <RANKING place="3" resultid="409" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6" agemax="21" agemin="18" name="Junioren weiblich">
                  <RANKINGS>
                    <RANKING place="2" resultid="44" />
                    <RANKING place="1" resultid="192" />
                    <RANKING place="3" resultid="385" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7" agemax="25" agemin="22" name="Pre-Master weiblich" />
                <AGEGROUP agegroupid="8" agemax="-1" agemin="26" name="Master weiblich">
                  <RANKINGS>
                    <RANKING place="1" resultid="112" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9" agemax="9" agemin="9" name="Kategorie E männlich" />
                <AGEGROUP agegroupid="10" agemax="11" agemin="10" name="Kategorie D männlich">
                  <RANKINGS>
                    <RANKING place="1" resultid="254" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11" agemax="13" agemin="12" name="Kategorie C männlich">
                  <RANKINGS>
                    <RANKING place="6" resultid="129" />
                    <RANKING place="5" resultid="166" />
                    <RANKING place="4" resultid="343" />
                    <RANKING place="2" resultid="359" />
                    <RANKING place="1" resultid="595" />
                    <RANKING place="3" resultid="599" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="12" agemax="15" agemin="14" name="Kategorie B männlich">
                  <RANKINGS>
                    <RANKING place="1" resultid="231" />
                    <RANKING place="3" resultid="350" />
                    <RANKING place="2" resultid="592" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="13" agemax="17" agemin="16" name="Kategorie A männlich">
                  <RANKINGS>
                    <RANKING place="3" resultid="270" />
                    <RANKING place="2" resultid="380" />
                    <RANKING place="1" resultid="423" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="14" agemax="21" agemin="18" name="Junioren männlich">
                  <RANKINGS>
                    <RANKING place="2" resultid="58" />
                    <RANKING place="3" resultid="494" />
                    <RANKING place="1" resultid="517" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15" agemax="25" agemin="22" name="Pre-Master männlich">
                  <RANKINGS>
                    <RANKING place="1" resultid="540" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="16" agemax="-1" agemin="26" name="Master männlich">
                  <RANKINGS>
                    <RANKING place="1" resultid="122" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="17" agemax="9" agemin="9" name="Kategorie E weiblich - LM" />
                <AGEGROUP agegroupid="18" agemax="11" agemin="10" name="Kategorie D weiblich - LM" />
                <AGEGROUP agegroupid="19" agemax="13" agemin="12" name="Kategorie C weiblich - LM" />
                <AGEGROUP agegroupid="20" agemax="15" agemin="14" name="Kategorie B weiblich - LM" />
                <AGEGROUP agegroupid="21" agemax="17" agemin="16" name="Kategorie A weiblich - LM" />
                <AGEGROUP agegroupid="22" agemax="21" agemin="18" name="Junioren weiblich - LM" />
                <AGEGROUP agegroupid="23" agemax="25" agemin="22" name="Pre-Master weiblich - LM" />
                <AGEGROUP agegroupid="24" agemax="-1" agemin="26" name="Master weiblich - LM" />
                <AGEGROUP agegroupid="25" agemax="9" agemin="9" name="Kategorie E männlich - LM" />
                <AGEGROUP agegroupid="26" agemax="11" agemin="10" name="Kategorie D männlich - LM" />
                <AGEGROUP agegroupid="27" agemax="13" agemin="12" name="Kategorie C männlich - LM" />
                <AGEGROUP agegroupid="28" agemax="15" agemin="14" name="Kategorie B männlich - LM" />
                <AGEGROUP agegroupid="29" agemax="17" agemin="16" name="Kategorie A männlich - LM">
                  <RANKINGS>
                    <RANKING place="1" resultid="270" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="30" agemax="21" agemin="18" name="Junioren männlich - LM">
                  <RANKINGS>
                    <RANKING place="2" resultid="494" />
                    <RANKING place="1" resultid="517" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="31" agemax="25" agemin="22" name="Pre-Master männlich - LM" />
                <AGEGROUP agegroupid="32" agemax="-1" agemin="26" name="Master männlich - LM" />
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="13" number="9" gender="X" round="TIM">
              <SWIMSTYLE stroke="SURFACE" relaycount="1" distance="200" />
              <FEE value="500" currency="EUR" />
              <HEATS>
                <HEAT heatid="13001" number="1" />
                <HEAT heatid="13002" number="2" />
                <HEAT heatid="13003" number="3" />
                <HEAT heatid="13004" number="4" />
                <HEAT heatid="13005" number="5" />
                <HEAT heatid="13006" number="6" />
                <HEAT heatid="13007" number="7" />
                <HEAT heatid="13008" number="8" />
                <HEAT heatid="13009" number="9" />
                <HEAT heatid="13010" number="10" />
                <HEAT heatid="13011" number="11" />
                <HEAT heatid="13012" number="12" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="9" agemin="9" name="Kategorie E weiblich">
                  <RANKINGS>
                    <RANKING place="3" resultid="54" />
                    <RANKING place="4" resultid="151" />
                    <RANKING place="5" resultid="217" />
                    <RANKING place="1" resultid="390" />
                    <RANKING place="2" resultid="461" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2" agemax="11" agemin="10" name="Kategorie D weiblich">
                  <RANKINGS>
                    <RANKING place="4" resultid="85" />
                    <RANKING place="16" resultid="143" />
                    <RANKING place="2" resultid="156" />
                    <RANKING place="6" resultid="172" />
                    <RANKING place="12" resultid="183" />
                    <RANKING place="10" resultid="188" />
                    <RANKING place="14" resultid="397" />
                    <RANKING place="13" resultid="413" />
                    <RANKING place="9" resultid="418" />
                    <RANKING place="7" resultid="469" />
                    <RANKING place="11" resultid="490" />
                    <RANKING place="15" resultid="513" />
                    <RANKING place="3" resultid="625" />
                    <RANKING place="5" resultid="629" />
                    <RANKING place="1" resultid="637" />
                    <RANKING place="8" resultid="649" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3" agemax="13" agemin="12" name="Kategorie C weiblich">
                  <RANKINGS>
                    <RANKING place="1" resultid="25" />
                    <RANKING place="2" resultid="65" />
                    <RANKING place="7" resultid="69" />
                    <RANKING place="3" resultid="73" />
                    <RANKING place="6" resultid="203" />
                    <RANKING place="4" resultid="235" />
                    <RANKING place="11" resultid="240" />
                    <RANKING place="8" resultid="266" />
                    <RANKING place="5" resultid="482" />
                    <RANKING place="10" resultid="577" />
                    <RANKING place="9" resultid="608" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="15" agemin="14" name="Kategorie B weiblich">
                  <RANKINGS>
                    <RANKING place="3" resultid="36" />
                    <RANKING place="1" resultid="504" />
                    <RANKING place="4" resultid="550" />
                    <RANKING place="2" resultid="569" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="17" agemin="16" name="Kategorie A weiblich">
                  <RANKINGS>
                    <RANKING place="5" resultid="91" />
                    <RANKING place="3" resultid="299" />
                    <RANKING place="2" resultid="426" />
                    <RANKING place="4" resultid="445" />
                    <RANKING place="6" resultid="581" />
                    <RANKING place="1" resultid="652" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6" agemax="21" agemin="18" name="Junioren weiblich">
                  <RANKINGS>
                    <RANKING place="4" resultid="5" />
                    <RANKING place="1" resultid="17" />
                    <RANKING place="2" resultid="62" />
                    <RANKING place="3" resultid="80" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7" agemax="25" agemin="22" name="Pre-Master weiblich" />
                <AGEGROUP agegroupid="8" agemax="-1" agemin="26" name="Master weiblich">
                  <RANKINGS>
                    <RANKING place="1" resultid="10" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9" agemax="9" agemin="9" name="Kategorie E männlich">
                  <RANKINGS>
                    <RANKING place="2" resultid="249" />
                    <RANKING place="3" resultid="372" />
                    <RANKING place="1" resultid="440" />
                    <RANKING place="4" resultid="465" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10" agemax="11" agemin="10" name="Kategorie D männlich">
                  <RANKINGS>
                    <RANKING place="4" resultid="330" />
                    <RANKING place="3" resultid="449" />
                    <RANKING place="2" resultid="457" />
                    <RANKING place="1" resultid="522" />
                    <RANKING place="5" resultid="544" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11" agemax="13" agemin="12" name="Kategorie C männlich">
                  <RANKINGS>
                    <RANKING place="8" resultid="31" />
                    <RANKING place="10" resultid="130" />
                    <RANKING place="9" resultid="167" />
                    <RANKING place="4" resultid="285" />
                    <RANKING place="7" resultid="326" />
                    <RANKING place="3" resultid="360" />
                    <RANKING place="5" resultid="436" />
                    <RANKING place="1" resultid="596" />
                    <RANKING place="2" resultid="600" />
                    <RANKING place="6" resultid="617" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="12" agemax="15" agemin="14" name="Kategorie B männlich">
                  <RANKINGS>
                    <RANKING place="4" resultid="40" />
                    <RANKING place="8" resultid="47" />
                    <RANKING place="9" resultid="76" />
                    <RANKING place="5" resultid="207" />
                    <RANKING place="2" resultid="278" />
                    <RANKING place="6" resultid="321" />
                    <RANKING place="1" resultid="474" />
                    <RANKING place="3" resultid="509" />
                    <RANKING place="7" resultid="535" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="13" agemax="17" agemin="16" name="Kategorie A männlich">
                  <RANKINGS>
                    <RANKING place="1" resultid="555" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="14" agemax="21" agemin="18" name="Junioren männlich">
                  <RANKINGS>
                    <RANKING place="1" resultid="486" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15" agemax="25" agemin="22" name="Pre-Master männlich">
                  <RANKINGS>
                    <RANKING place="1" resultid="317" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="16" agemax="-1" agemin="26" name="Master männlich" />
                <AGEGROUP agegroupid="17" agemax="9" agemin="9" name="Kategorie E weiblich - LM">
                  <RANKINGS>
                    <RANKING place="1" resultid="461" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="18" agemax="11" agemin="10" name="Kategorie D weiblich - LM">
                  <RANKINGS>
                    <RANKING place="1" resultid="469" />
                    <RANKING place="2" resultid="490" />
                    <RANKING place="3" resultid="513" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="19" agemax="13" agemin="12" name="Kategorie C weiblich - LM">
                  <RANKINGS>
                    <RANKING place="2" resultid="266" />
                    <RANKING place="1" resultid="482" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="20" agemax="15" agemin="14" name="Kategorie B weiblich - LM">
                  <RANKINGS>
                    <RANKING place="1" resultid="504" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="21" agemax="17" agemin="16" name="Kategorie A weiblich - LM">
                  <RANKINGS>
                    <RANKING place="2" resultid="299" />
                    <RANKING place="3" resultid="445" />
                    <RANKING place="1" resultid="652" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="22" agemax="21" agemin="18" name="Junioren weiblich - LM" />
                <AGEGROUP agegroupid="23" agemax="25" agemin="22" name="Pre-Master weiblich - LM" />
                <AGEGROUP agegroupid="24" agemax="-1" agemin="26" name="Master weiblich - LM" />
                <AGEGROUP agegroupid="25" agemax="9" agemin="9" name="Kategorie E männlich - LM">
                  <RANKINGS>
                    <RANKING place="1" resultid="440" />
                    <RANKING place="2" resultid="465" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="26" agemax="11" agemin="10" name="Kategorie D männlich - LM">
                  <RANKINGS>
                    <RANKING place="4" resultid="330" />
                    <RANKING place="3" resultid="449" />
                    <RANKING place="2" resultid="457" />
                    <RANKING place="1" resultid="522" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="27" agemax="13" agemin="12" name="Kategorie C männlich - LM">
                  <RANKINGS>
                    <RANKING place="1" resultid="285" />
                    <RANKING place="3" resultid="326" />
                    <RANKING place="2" resultid="436" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="28" agemax="15" agemin="14" name="Kategorie B männlich - LM">
                  <RANKINGS>
                    <RANKING place="2" resultid="278" />
                    <RANKING place="4" resultid="321" />
                    <RANKING place="1" resultid="474" />
                    <RANKING place="3" resultid="509" />
                    <RANKING place="5" resultid="535" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="29" agemax="17" agemin="16" name="Kategorie A männlich - LM" />
                <AGEGROUP agegroupid="30" agemax="21" agemin="18" name="Junioren männlich - LM">
                  <RANKINGS>
                    <RANKING place="1" resultid="486" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="31" agemax="25" agemin="22" name="Pre-Master männlich - LM">
                  <RANKINGS>
                    <RANKING place="1" resultid="317" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="32" agemax="-1" agemin="26" name="Master männlich - LM" />
                <AGEGROUP agegroupid="33" agemax="8" agemin="0" name="Jg. 2015 u. jünger">
                  <RANKINGS>
                    <RANKING place="2" resultid="257" />
                    <RANKING place="3" resultid="639" />
                    <RANKING place="1" resultid="645" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="14" number="10" gender="X" round="TIM">
              <SWIMSTYLE stroke="UNKNOWN" relaycount="4" distance="100" />
              <FEE value="750" currency="EUR" />
              <HEATS>
                <HEAT heatid="14001" number="1" />
                <HEAT heatid="14002" number="2" />
                <HEAT heatid="14003" number="3" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="3" agemax="14" agemin="0" name="Kategorie C">
                  <RANKINGS>
                    <RANKING place="2" resultid="19" />
                    <RANKING place="7" resultid="209" />
                    <RANKING place="5" resultid="364" />
                    <RANKING place="6" resultid="365" />
                    <RANKING place="1" resultid="559" />
                    <RANKING place="3" resultid="560" />
                    <RANKING place="4" resultid="561" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2" agemax="19" agemin="15" name="Kategorie B">
                  <RANKINGS>
                    <RANKING place="1" resultid="18" />
                    <RANKING place="5" resultid="20" />
                    <RANKING place="7" resultid="21" />
                    <RANKING place="3" resultid="208" />
                    <RANKING place="4" resultid="259" />
                    <RANKING place="6" resultid="366" />
                    <RANKING place="9" resultid="367" />
                    <RANKING place="8" resultid="368" />
                    <RANKING place="2" resultid="536" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1" agemax="-1" agemin="20" name="Kategorie A">
                  <RANKINGS>
                    <RANKING place="2" resultid="92" />
                    <RANKING place="1" resultid="258" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
          </EVENTS>
        </SESSION>
      </SESSIONS>
      <CLUBS>
        <CLUB name="1. Chemnitzer Tauchverein e.V." nation="GER" region="20" code="0">
          <ATHLETES>
            <ATHLETE athleteid="132" birthdate="2006-01-01" gender="M" lastname="Lorenz" firstname="Emil" license="0">
              <RESULTS>
                <RESULT resultid="420" eventid="1" swimtime="00:00:16.51" lane="6" heatid="1007" />
                <RESULT resultid="421" eventid="5" swimtime="00:00:42.08" lane="6" heatid="5018" />
                <RESULT resultid="422" eventid="10" swimtime="00:00:18.94" lane="7" heatid="10018" />
                <RESULT resultid="423" eventid="12" swimtime="00:00:42.71" lane="6" heatid="12005" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="133" birthdate="2007-01-01" gender="F" lastname="Ullrich" firstname="Johanna Hermine" license="0">
              <RESULTS>
                <RESULT resultid="424" eventid="3" swimtime="00:04:05.05" lane="1" heatid="3009">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:54.50" />
                    <SPLIT distance="200" swimtime="00:01:58.92" />
                    <SPLIT distance="300" swimtime="00:03:03.90" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="425" eventid="5" status="DSQ" swimtime="00:00:53.60" lane="2" heatid="5014" comment="falscher Start" />
                <RESULT resultid="426" eventid="13" swimtime="00:01:55.29" lane="2" heatid="13010">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:55.26" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="134" birthdate="1997-01-01" gender="F" lastname="Brinster" firstname="Luise" license="0">
              <RESULTS>
                <RESULT resultid="427" eventid="3" swimtime="00:04:38.69" lane="3" heatid="3008">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:03.10" />
                    <SPLIT distance="200" swimtime="00:02:14.67" />
                    <SPLIT distance="300" swimtime="00:03:27.69" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="428" eventid="10" swimtime="00:00:26.07" lane="8" heatid="10012" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="135" birthdate="2005-01-01" gender="M" lastname="Porges" firstname="Marcel" license="0">
              <RESULTS>
                <RESULT resultid="429" eventid="1" swimtime="00:00:16.14" lane="5" heatid="1007" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="136" birthdate="1998-01-01" gender="F" lastname="Oehme" firstname="Victoria" license="0">
              <RESULTS>
                <RESULT resultid="430" eventid="1" status="DNS" swimtime="00:00:00.00" lane="4" heatid="1001" />
                <RESULT resultid="431" eventid="5" swimtime="00:00:57.95" lane="4" heatid="5011" />
                <RESULT resultid="432" eventid="10" status="DNS" swimtime="00:00:00.00" lane="7" heatid="10010" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY number="1" gender="X" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="419" eventid="14" status="DSQ" swimtime="00:02:33.73" lane="2" heatid="14001" comment="Falscher Start.">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:51.20" />
                    <SPLIT distance="200" swimtime="00:01:47.68" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="136" number="1" />
                    <RELAYPOSITION athleteid="134" number="2" />
                    <RELAYPOSITION athleteid="133" number="3" />
                    <RELAYPOSITION athleteid="132" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB name="Binger Tauchsportclub e.V." nation="GER" region="29" code="0">
          <ATHLETES>
            <ATHLETE athleteid="1" birthdate="2004-01-01" gender="F" lastname="Walter" firstname="Julia" license="0">
              <RESULTS>
                <RESULT resultid="1" eventid="1" swimtime="00:00:23.09" lane="5" heatid="1003" />
                <RESULT resultid="2" eventid="3" swimtime="00:04:16.38" lane="4" heatid="3009">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:57.91" />
                    <SPLIT distance="200" swimtime="00:02:02.76" />
                    <SPLIT distance="300" swimtime="00:03:09.17" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="3" eventid="5" swimtime="00:00:54.98" lane="4" heatid="5015" />
                <RESULT resultid="4" eventid="10" status="DSQ" swimtime="00:00:24.82" lane="6" heatid="10014" comment="falscher Start" />
                <RESULT resultid="5" eventid="13" swimtime="00:02:02.25" lane="4" heatid="13011">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:57.62" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="2" birthdate="1997-01-01" gender="F" lastname="Walter" firstname="Lisa" license="0">
              <RESULTS>
                <RESULT resultid="6" eventid="1" swimtime="00:00:24.55" lane="3" heatid="1002" />
                <RESULT resultid="7" eventid="3" swimtime="00:04:22.16" lane="4" heatid="3008">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:00.93" />
                    <SPLIT distance="200" swimtime="00:02:06.97" />
                    <SPLIT distance="300" swimtime="00:03:15.00" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="8" eventid="5" swimtime="00:00:56.00" lane="1" heatid="5014" />
                <RESULT resultid="9" eventid="10" swimtime="00:00:25.42" lane="4" heatid="10012" />
                <RESULT resultid="10" eventid="13" swimtime="00:02:03.57" lane="1" heatid="13011">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:00.21" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="SC DHfK Leipzig Flossenschwimmen" nation="GER" region="20" code="0">
          <ATHLETES>
            <ATHLETE athleteid="3" birthdate="2001-01-01" gender="F" lastname="Hecke" firstname="Aimee Joy" license="0">
              <RESULTS>
                <RESULT resultid="11" eventid="5" swimtime="00:00:45.32" lane="5" heatid="5016" />
                <RESULT resultid="12" eventid="10" swimtime="00:00:20.69" lane="3" heatid="10017" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="4" birthdate="2003-01-01" gender="F" lastname="Fischer" firstname="Josefine" license="0">
              <RESULTS>
                <RESULT resultid="13" eventid="1" swimtime="00:00:20.49" lane="8" heatid="1004" />
                <RESULT resultid="14" eventid="10" swimtime="00:00:21.51" lane="7" heatid="10015" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="5" birthdate="2004-01-01" gender="F" lastname="Barthel" firstname="Nadja" license="0">
              <RESULTS>
                <RESULT resultid="15" eventid="5" swimtime="00:00:41.50" lane="3" heatid="5018" />
                <RESULT resultid="16" eventid="10" status="DSQ" swimtime="00:00:19.05" lane="6" heatid="10018" comment="Tauchzüge außerhalb der 15m-Zone" />
                <RESULT resultid="17" eventid="13" swimtime="00:01:35.23" lane="4" heatid="13012">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:46.50" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="SSC Halle" nation="GER" region="27" code="0">
          <ATHLETES>
            <ATHLETE athleteid="80" birthdate="2012-01-01" gender="M" lastname="Anacker" firstname="Caylan" license="0">
              <RESULTS>
                <RESULT resultid="261" eventid="5" swimtime="00:01:39.04" lane="3" heatid="5001" />
                <RESULT resultid="262" eventid="8" swimtime="00:00:49.27" lane="5" heatid="8001" />
                <RESULT resultid="263" eventid="10" swimtime="00:00:42.41" lane="3" heatid="10001" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="81" birthdate="2011-01-01" gender="F" lastname="Richter" firstname="Charlotte" license="0">
              <RESULTS>
                <RESULT resultid="264" eventid="5" swimtime="00:01:14.79" lane="8" heatid="5004" />
                <RESULT resultid="265" eventid="10" status="DSQ" swimtime="00:00:32.39" lane="4" heatid="10003" comment="falscher Start" />
                <RESULT resultid="266" eventid="13" swimtime="00:02:52.93" lane="1" heatid="13004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:25.80" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="82" birthdate="2007-01-01" gender="M" lastname="Koch" firstname="Elias" license="0">
              <RESULTS>
                <RESULT resultid="267" eventid="1" swimtime="00:00:19.38" lane="2" heatid="1006" />
                <RESULT resultid="268" eventid="5" swimtime="00:00:48.92" lane="1" heatid="5017" />
                <RESULT resultid="269" eventid="10" swimtime="00:00:21.29" lane="7" heatid="10017" />
                <RESULT resultid="270" eventid="12" swimtime="00:00:50.65" lane="6" heatid="12004" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="83" birthdate="2015-01-01" gender="M" lastname="Streblow" firstname="Emil" license="0">
              <RESULTS>
                <RESULT resultid="271" eventid="2" swimtime="00:00:49.94" lane="6" heatid="2001" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="84" birthdate="2010-01-01" gender="M" lastname="Eichberg" firstname="Eric" license="0">
              <RESULTS>
                <RESULT resultid="272" eventid="5" status="DNS" swimtime="00:00:00.00" lane="1" heatid="5006" />
                <RESULT resultid="273" eventid="10" status="DNS" swimtime="00:00:00.00" lane="5" heatid="10006" />
                <RESULT resultid="274" eventid="13" status="DNS" swimtime="00:00:00.00" lane="8" heatid="13007" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="85" birthdate="2008-01-01" gender="M" lastname="Baumbach" firstname="Felix" license="0">
              <RESULTS>
                <RESULT resultid="275" eventid="3" swimtime="00:04:09.83" lane="2" heatid="3009">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:57.72" />
                    <SPLIT distance="200" swimtime="00:02:02.25" />
                    <SPLIT distance="300" swimtime="00:03:08.13" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="276" eventid="5" swimtime="00:00:52.10" lane="2" heatid="5015" />
                <RESULT resultid="277" eventid="10" swimtime="00:00:23.21" lane="5" heatid="10015" />
                <RESULT resultid="278" eventid="13" swimtime="00:01:54.71" lane="7" heatid="13011">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:55.12" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="86" birthdate="2013-01-01" gender="M" lastname="Rosemann" firstname="Henri" license="0">
              <RESULTS>
                <RESULT resultid="279" eventid="5" status="DSQ" swimtime="00:01:15.05" lane="6" heatid="5006" comment="Falscher Start." />
                <RESULT resultid="280" eventid="8" swimtime="00:00:44.98" lane="1" heatid="8004" />
                <RESULT resultid="281" eventid="10" swimtime="00:00:36.00" lane="3" heatid="10003" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="87" birthdate="2011-01-01" gender="M" lastname="Reinicke" firstname="Jakob" license="0">
              <RESULTS>
                <RESULT resultid="282" eventid="3" swimtime="00:05:15.19" lane="8" heatid="3006">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:12.73" />
                    <SPLIT distance="200" swimtime="00:02:33.94" />
                    <SPLIT distance="300" swimtime="00:03:56.29" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="283" eventid="5" swimtime="00:01:00.23" lane="1" heatid="5012" />
                <RESULT resultid="284" eventid="10" swimtime="00:00:25.74" lane="5" heatid="10011" />
                <RESULT resultid="285" eventid="13" swimtime="00:02:14.59" lane="1" heatid="13009">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:05.08" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="88" birthdate="2016-01-01" gender="M" lastname="Gernhardt" firstname="Justus" license="0">
              <RESULTS>
                <RESULT resultid="286" eventid="2" swimtime="00:01:13.84" lane="3" heatid="2001" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="89" birthdate="2010-01-01" gender="M" lastname="Harms" firstname="Justus" license="0">
              <RESULTS>
                <RESULT resultid="287" eventid="3" status="DNS" swimtime="00:00:00.00" lane="5" heatid="3005" />
                <RESULT resultid="288" eventid="5" status="DNS" swimtime="00:00:00.00" lane="5" heatid="5011" />
                <RESULT resultid="289" eventid="10" status="DNS" swimtime="00:00:00.00" lane="2" heatid="10010" />
                <RESULT resultid="290" eventid="13" status="DNS" swimtime="00:00:00.00" lane="5" heatid="13007" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="90" birthdate="2014-01-01" gender="F" lastname="Friess" firstname="Klara" license="0">
              <RESULTS>
                <RESULT resultid="291" eventid="5" status="DNS" swimtime="00:00:00.00" lane="8" heatid="5002" />
                <RESULT resultid="292" eventid="8" status="DNS" swimtime="00:00:00.00" lane="8" heatid="8002" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="91" birthdate="2007-01-01" gender="F" lastname="Gallitz" firstname="Laura" license="0">
              <RESULTS>
                <RESULT resultid="293" eventid="1" status="DSQ" swimtime="00:00:26.41" lane="1" heatid="1003" comment="Aufgabe nach 35 m (aufgetaucht)" />
                <RESULT resultid="294" eventid="5" swimtime="00:00:57.54" lane="2" heatid="5012" />
                <RESULT resultid="295" eventid="10" swimtime="00:00:24.81" lane="6" heatid="10013" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="92" birthdate="2006-01-01" gender="F" lastname="Dietrich" firstname="Lea" license="0">
              <RESULTS>
                <RESULT resultid="296" eventid="1" swimtime="00:00:19.46" lane="4" heatid="1005" />
                <RESULT resultid="297" eventid="5" swimtime="00:00:48.22" lane="4" heatid="5016" />
                <RESULT resultid="298" eventid="10" swimtime="00:00:21.90" lane="1" heatid="10017" />
                <RESULT resultid="299" eventid="13" swimtime="00:01:56.97" lane="2" heatid="13012">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:54.05" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="93" birthdate="2014-01-01" gender="F" lastname="Keck" firstname="Lilly" license="0">
              <RESULTS>
                <RESULT resultid="300" eventid="5" status="DSQ" swimtime="00:00:00.00" lane="1" heatid="5002" comment="Falscher Start.&#xA;Aufgabe bei 50m." />
                <RESULT resultid="301" eventid="8" swimtime="00:00:43.57" lane="4" heatid="8001" />
                <RESULT resultid="302" eventid="10" swimtime="00:00:38.19" lane="5" heatid="10001" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="94" birthdate="2016-01-01" gender="M" lastname="Krüger" firstname="Matheo" license="0">
              <RESULTS>
                <RESULT resultid="303" eventid="2" swimtime="00:01:13.43" lane="4" heatid="2001" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="95" birthdate="2013-01-01" gender="F" lastname="Stephan" firstname="Mathilda" license="0">
              <RESULTS>
                <RESULT resultid="304" eventid="5" swimtime="00:01:38.08" lane="4" heatid="5002" />
                <RESULT resultid="305" eventid="8" swimtime="00:00:51.52" lane="1" heatid="8002" />
                <RESULT resultid="306" eventid="10" swimtime="00:00:43.13" lane="7" heatid="10002" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="96" birthdate="2000-01-01" gender="M" lastname="Kubler" firstname="Max" license="0">
              <RESULTS>
                <RESULT resultid="307" eventid="1" swimtime="00:00:18.38" lane="3" heatid="1005" />
                <RESULT resultid="308" eventid="5" swimtime="00:00:47.84" lane="7" heatid="5015" />
                <RESULT resultid="309" eventid="10" swimtime="00:00:22.00" lane="2" heatid="10015" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="97" birthdate="2014-01-01" gender="M" lastname="Frenzel" firstname="Nick" license="0">
              <RESULTS>
                <RESULT resultid="310" eventid="5" status="DSQ" swimtime="00:01:31.05" lane="4" heatid="5003" comment="Falsche Ausrüstung (kein Schnorchel)" />
                <RESULT resultid="311" eventid="8" status="DSQ" swimtime="00:00:46.38" lane="2" heatid="8002" comment="falscher Schwimmstil - mehrere Wechselbeinschläge nach dem Start" />
                <RESULT resultid="312" eventid="10" swimtime="00:00:40.09" lane="2" heatid="10002" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="98" birthdate="2015-01-01" gender="M" lastname="Kathmann" firstname="Niels" license="0">
              <RESULTS>
                <RESULT resultid="313" eventid="2" swimtime="00:00:52.29" lane="5" heatid="2001" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="99" birthdate="2001-01-01" gender="M" lastname="Heidari" firstname="Parsa" license="0">
              <RESULTS>
                <RESULT resultid="314" eventid="1" status="DSQ" swimtime="00:00:00.00" lane="1" heatid="1005" comment="falscher Start" />
                <RESULT resultid="315" eventid="5" swimtime="00:00:49.01" lane="7" heatid="5016" />
                <RESULT resultid="316" eventid="10" swimtime="00:00:22.42" lane="2" heatid="10016" />
                <RESULT resultid="317" eventid="13" swimtime="00:01:48.58" lane="6" heatid="13011">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:51.11" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="100" birthdate="2009-01-01" gender="M" lastname="Gaudig" firstname="Paul" license="0">
              <RESULTS>
                <RESULT resultid="318" eventid="1" swimtime="00:00:22.95" lane="3" heatid="1003" />
                <RESULT resultid="319" eventid="5" swimtime="00:00:56.54" lane="8" heatid="5014" />
                <RESULT resultid="320" eventid="10" swimtime="00:00:23.62" lane="6" heatid="10015" />
                <RESULT resultid="321" eventid="13" swimtime="00:02:13.69" lane="1" heatid="13010">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:01.89" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="101" birthdate="2003-01-01" gender="M" lastname="Gerlach" firstname="Ruben" license="0">
              <RESULTS>
                <RESULT resultid="322" eventid="1" swimtime="00:00:18.37" lane="1" heatid="1006" />
                <RESULT resultid="323" eventid="10" swimtime="00:00:20.37" lane="5" heatid="10017" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="102" birthdate="2011-01-01" gender="M" lastname="Frenzel" firstname="Tim" license="0">
              <RESULTS>
                <RESULT resultid="324" eventid="5" swimtime="00:01:10.21" lane="2" heatid="5008" />
                <RESULT resultid="325" eventid="10" status="DSQ" swimtime="00:00:30.36" lane="4" heatid="10008" comment="falscher Start" />
                <RESULT resultid="326" eventid="13" swimtime="00:02:29.29" lane="5" heatid="13006">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:14.43" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="103" birthdate="2012-01-01" gender="M" lastname="Gaudig" firstname="Tom" license="0">
              <RESULTS>
                <RESULT resultid="327" eventid="5" swimtime="00:01:12.06" lane="1" heatid="5008" />
                <RESULT resultid="328" eventid="8" swimtime="00:00:35.08" lane="1" heatid="8003" />
                <RESULT resultid="329" eventid="10" swimtime="00:00:31.92" lane="8" heatid="10005" />
                <RESULT resultid="330" eventid="13" swimtime="00:02:44.29" lane="3" heatid="13005">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:22.76" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="192" birthdate="2007-01-01" gender="F" lastname="Gerlach" firstname="Meret" license="0">
              <RESULTS>
                <RESULT resultid="651" eventid="1" swimtime="00:00:21.07" lane="4" heatid="1004" />
                <RESULT resultid="652" eventid="13" swimtime="00:01:48.69" lane="7" heatid="13012">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:52.50" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY number="1" gender="X" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="258" eventid="14" swimtime="00:02:20.93" lane="3" heatid="14003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:44.71" />
                    <SPLIT distance="200" swimtime="00:01:33.92" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="99" number="1" />
                    <RELAYPOSITION athleteid="92" number="2" />
                    <RELAYPOSITION athleteid="82" number="3" />
                    <RELAYPOSITION athleteid="192" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="2" gender="X" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="259" eventid="14" swimtime="00:02:49.12" lane="2" heatid="14003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:49.85" />
                    <SPLIT distance="200" swimtime="00:01:46.42" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="91" number="1" />
                    <RELAYPOSITION athleteid="85" number="2" />
                    <RELAYPOSITION athleteid="100" number="3" />
                    <RELAYPOSITION athleteid="81" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="3" gender="X" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="260" eventid="14" status="DNS" swimtime="00:00:00.00" lane="7" heatid="14002">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="89" number="1" />
                    <RELAYPOSITION athleteid="87" number="2" />
                    <RELAYPOSITION athleteid="102" number="3" />
                    <RELAYPOSITION athleteid="86" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB name="Startgemeinschaft Dresden" nation="GER" region="20" code="0">
          <ATHLETES>
            <ATHLETE athleteid="29" birthdate="2013-01-01" gender="F" lastname="Stegemann" firstname="Anna" license="0">
              <RESULTS>
                <RESULT resultid="93" eventid="5" swimtime="00:01:14.99" lane="2" heatid="5004" />
                <RESULT resultid="94" eventid="10" status="DSQ" swimtime="00:00:32.18" lane="4" heatid="10002" comment="falscher Start" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="30" birthdate="2009-01-01" gender="M" lastname="Hübner" firstname="Christoph" license="0">
              <RESULTS>
                <RESULT resultid="95" eventid="5" swimtime="00:01:18.03" lane="2" heatid="5006" />
                <RESULT resultid="96" eventid="10" status="DSQ" swimtime="00:00:29.28" lane="4" heatid="10006" comment="falscher Start" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="31" birthdate="2010-01-01" gender="F" lastname="Reichel" firstname="Emily" license="0">
              <RESULTS>
                <RESULT resultid="97" eventid="5" status="DNS" swimtime="00:00:00.00" lane="2" heatid="5010" />
                <RESULT resultid="98" eventid="10" status="DNS" swimtime="00:00:00.00" lane="8" heatid="10010" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="32" birthdate="2010-01-01" gender="F" lastname="Mucha" firstname="Helene" license="0">
              <RESULTS>
                <RESULT resultid="99" eventid="5" swimtime="00:01:11.58" lane="5" heatid="5005" />
                <RESULT resultid="100" eventid="10" swimtime="00:00:32.09" lane="3" heatid="10005" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="33" birthdate="2006-01-01" gender="F" lastname="Schürer" firstname="Katka" license="0">
              <RESULTS>
                <RESULT resultid="101" eventid="5" swimtime="00:01:07.61" lane="5" heatid="5008" />
                <RESULT resultid="102" eventid="10" swimtime="00:00:30.68" lane="4" heatid="10007" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="34" birthdate="2007-01-01" gender="F" lastname="Marquardt" firstname="Lotte" license="0">
              <RESULTS>
                <RESULT resultid="103" eventid="1" swimtime="00:00:25.30" lane="2" heatid="1002" />
                <RESULT resultid="104" eventid="5" swimtime="00:00:59.61" lane="7" heatid="5011" />
                <RESULT resultid="105" eventid="10" swimtime="00:00:27.37" lane="5" heatid="10010" />
                <RESULT resultid="106" eventid="12" swimtime="00:01:00.58" lane="2" heatid="12002" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="35" birthdate="2011-01-01" gender="M" lastname="Buchmann" firstname="Marco" license="0">
              <RESULTS>
                <RESULT resultid="107" eventid="5" swimtime="00:01:11.84" lane="4" heatid="5006" />
                <RESULT resultid="108" eventid="10" swimtime="00:00:31.41" lane="8" heatid="10006" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="36" birthdate="1986-01-01" gender="F" lastname="Klar" firstname="Margarethe" license="0">
              <RESULTS>
                <RESULT resultid="109" eventid="3" swimtime="00:04:46.84" lane="3" heatid="3007">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:04.90" />
                    <SPLIT distance="200" swimtime="00:02:18.79" />
                    <SPLIT distance="300" swimtime="00:03:34.65" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="110" eventid="6" swimtime="00:04:42.51" lane="2" heatid="6001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:04.10" />
                    <SPLIT distance="200" swimtime="00:02:16.14" />
                    <SPLIT distance="300" swimtime="00:03:32.12" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="111" eventid="10" swimtime="00:00:30.42" lane="3" heatid="10010" />
                <RESULT resultid="112" eventid="12" swimtime="00:01:01.86" lane="6" heatid="12003" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="37" birthdate="2011-01-01" gender="F" lastname="Oehme" firstname="Mia" license="0">
              <RESULTS>
                <RESULT resultid="113" eventid="5" swimtime="00:01:11.79" lane="3" heatid="5008" />
                <RESULT resultid="114" eventid="10" swimtime="00:00:32.08" lane="8" heatid="10007" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="38" birthdate="2011-01-01" gender="F" lastname="Müller" firstname="Reni" license="0">
              <RESULTS>
                <RESULT resultid="115" eventid="5" swimtime="00:01:08.49" lane="7" heatid="5007" />
                <RESULT resultid="116" eventid="10" swimtime="00:00:32.17" lane="3" heatid="10007" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="39" birthdate="2007-01-01" gender="F" lastname="Razumovska" firstname="Sophiya" license="0">
              <RESULTS>
                <RESULT resultid="117" eventid="1" status="DSQ" swimtime="00:00:24.85" lane="3" heatid="1001" comment="falscher Start" />
                <RESULT resultid="118" eventid="5" swimtime="00:01:04.71" lane="7" heatid="5010" />
                <RESULT resultid="119" eventid="10" swimtime="00:00:27.20" lane="3" heatid="10009" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="40" birthdate="1978-01-01" gender="M" lastname="Hoffmann" firstname="Stefan" license="0">
              <RESULTS>
                <RESULT resultid="120" eventid="1" swimtime="00:00:19.17" lane="8" heatid="1006" />
                <RESULT resultid="121" eventid="10" swimtime="00:00:22.88" lane="1" heatid="10015" />
                <RESULT resultid="122" eventid="12" swimtime="00:00:45.49" lane="3" heatid="12004" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY number="1" gender="X" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="92" eventid="14" swimtime="00:02:53.78" lane="5" heatid="14002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:47.81" />
                    <SPLIT distance="200" swimtime="00:01:51.42" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="40" number="1" />
                    <RELAYPOSITION athleteid="34" number="2" />
                    <RELAYPOSITION athleteid="36" number="3" />
                    <RELAYPOSITION athleteid="39" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB name="Tauchclub NEMO Plauen e.V." nation="GER" region="20" code="0">
          <ATHLETES>
            <ATHLETE athleteid="188" birthdate="2009-01-01" gender="F" lastname="Troppschuh" firstname="Hannah" license="0">
              <RESULTS>
                <RESULT resultid="630" eventid="1" swimtime="00:00:19.72" lane="3" heatid="1006" />
                <RESULT resultid="631" eventid="5" swimtime="00:00:47.19" lane="3" heatid="5017" />
                <RESULT resultid="632" eventid="10" swimtime="00:00:22.63" lane="8" heatid="10017" />
                <RESULT resultid="633" eventid="12" swimtime="00:00:47.87" lane="2" heatid="12005" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="189" birthdate="2012-01-01" gender="F" lastname="Troppschuh" firstname="Lotte" license="0">
              <RESULTS>
                <RESULT resultid="634" eventid="5" swimtime="00:00:50.55" lane="4" heatid="5014" />
                <RESULT resultid="635" eventid="8" swimtime="00:00:26.33" lane="4" heatid="8004" />
                <RESULT resultid="636" eventid="10" swimtime="00:00:22.66" lane="4" heatid="10013" />
                <RESULT resultid="637" eventid="13" swimtime="00:02:04.43" lane="5" heatid="13009">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:00.01" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="Tauchsportclub Erfurt e.V." nation="GER" region="35" code="0">
          <ATHLETES>
            <ATHLETE athleteid="171" birthdate="2010-01-01" gender="F" lastname="Abe" firstname="Adina" license="0">
              <RESULTS>
                <RESULT resultid="562" eventid="3" swimtime="00:04:20.76" lane="6" heatid="3008">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:00.79" />
                    <SPLIT distance="200" swimtime="00:02:08.26" />
                    <SPLIT distance="300" swimtime="00:03:17.05" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="563" eventid="5" swimtime="00:00:53.85" lane="3" heatid="5015" />
                <RESULT resultid="564" eventid="10" status="DNS" swimtime="00:00:00.00" lane="7" heatid="10014" />
                <RESULT resultid="565" eventid="12" swimtime="00:00:52.12" lane="8" heatid="12004" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="172" birthdate="2009-01-01" gender="F" lastname="Darzhaniia" firstname="Alisa" license="0">
              <RESULTS>
                <RESULT resultid="566" eventid="3" swimtime="00:03:59.00" lane="5" heatid="3009">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:53.21" />
                    <SPLIT distance="200" swimtime="00:01:54.49" />
                    <SPLIT distance="300" swimtime="00:02:59.18" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="567" eventid="5" swimtime="00:00:49.59" lane="6" heatid="5016" />
                <RESULT resultid="568" eventid="10" swimtime="00:00:22.22" lane="5" heatid="10016" />
                <RESULT resultid="569" eventid="13" swimtime="00:01:52.35" lane="8" heatid="13012">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:53.07" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="173" birthdate="2009-01-01" gender="F" lastname="Zitzmann" firstname="Annalena" license="0">
              <RESULTS>
                <RESULT resultid="570" eventid="1" swimtime="00:00:21.60" lane="4" heatid="1003" />
                <RESULT resultid="571" eventid="3" status="DSQ" swimtime="00:04:22.18" lane="8" heatid="3007" comment="15 m nach Start übertaucht">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:59.32" />
                    <SPLIT distance="200" swimtime="00:02:07.60" />
                    <SPLIT distance="300" swimtime="00:03:17.32" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="572" eventid="5" swimtime="00:00:51.93" lane="6" heatid="5015" />
                <RESULT resultid="573" eventid="10" swimtime="00:00:22.54" lane="4" heatid="10015" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="174" birthdate="2010-01-01" gender="F" lastname="Hartung" firstname="Antonia Lea" license="0">
              <RESULTS>
                <RESULT resultid="574" eventid="3" swimtime="00:06:10.21" lane="5" heatid="3001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:23.68" />
                    <SPLIT distance="200" swimtime="00:03:01.45" />
                    <SPLIT distance="300" swimtime="00:04:40.74" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="575" eventid="5" swimtime="00:01:13.85" lane="3" heatid="5004" />
                <RESULT resultid="576" eventid="10" swimtime="00:00:32.60" lane="6" heatid="10004" />
                <RESULT resultid="577" eventid="13" swimtime="00:03:04.32" lane="7" heatid="13004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:26.93" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="175" birthdate="2007-01-01" gender="F" lastname="Zieger" firstname="Emilie" license="0">
              <RESULTS>
                <RESULT resultid="578" eventid="3" swimtime="00:05:01.87" lane="6" heatid="3005">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:08.15" />
                    <SPLIT distance="200" swimtime="00:02:27.76" />
                    <SPLIT distance="300" swimtime="00:03:48.67" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="579" eventid="5" status="DSQ" swimtime="00:01:06.91" lane="4" heatid="5010" comment="falscher Start" />
                <RESULT resultid="580" eventid="10" swimtime="00:00:32.11" lane="4" heatid="10009" />
                <RESULT resultid="581" eventid="13" swimtime="00:02:24.65" lane="2" heatid="13008">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:09.43" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="176" birthdate="2014-01-01" gender="F" lastname="Wagner" firstname="Emma" license="0">
              <RESULTS>
                <RESULT resultid="582" eventid="5" status="DNS" swimtime="00:00:00.00" lane="2" heatid="5001" />
                <RESULT resultid="583" eventid="8" status="DNS" swimtime="00:00:00.00" lane="1" heatid="8001" />
                <RESULT resultid="584" eventid="10" status="DNS" swimtime="00:00:00.00" lane="7" heatid="10001" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="177" birthdate="2009-01-01" gender="F" lastname="Henkel" firstname="Friederike" license="0">
              <RESULTS>
                <RESULT resultid="585" eventid="1" status="DSQ" swimtime="00:00:00.00" lane="6" heatid="1001" comment="Aufgegeben nach 35 m" />
                <RESULT resultid="586" eventid="3" swimtime="00:05:11.61" lane="1" heatid="3005">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:08.97" />
                    <SPLIT distance="200" swimtime="00:02:30.88" />
                    <SPLIT distance="300" swimtime="00:03:54.39" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="587" eventid="10" swimtime="00:00:26.30" lane="1" heatid="10012" />
                <RESULT resultid="588" eventid="12" swimtime="00:01:02.58" lane="4" heatid="12001" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="178" birthdate="2009-01-01" gender="M" lastname="Artschwager" firstname="Gustaf" license="0">
              <RESULTS>
                <RESULT resultid="589" eventid="1" swimtime="00:00:27.16" lane="2" heatid="1001" />
                <RESULT resultid="590" eventid="3" swimtime="00:04:41.75" lane="2" heatid="3006">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:05.41" />
                    <SPLIT distance="200" swimtime="00:02:19.05" />
                    <SPLIT distance="300" swimtime="00:03:33.79" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="591" eventid="10" swimtime="00:00:27.87" lane="4" heatid="10011" />
                <RESULT resultid="592" eventid="12" swimtime="00:01:11.25" lane="8" heatid="12002" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="179" birthdate="2010-01-01" gender="M" lastname="Leipold" firstname="Jakob" license="0">
              <RESULTS>
                <RESULT resultid="593" eventid="5" swimtime="00:00:53.72" lane="7" heatid="5014" />
                <RESULT resultid="594" eventid="10" swimtime="00:00:25.47" lane="8" heatid="10014" />
                <RESULT resultid="595" eventid="12" swimtime="00:00:52.61" lane="4" heatid="12003" />
                <RESULT resultid="596" eventid="13" swimtime="00:02:07.47" lane="3" heatid="13010">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:01.16" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="180" birthdate="2010-01-01" gender="M" lastname="Hochstein" firstname="Jean Paul" license="0">
              <RESULTS>
                <RESULT resultid="597" eventid="5" swimtime="00:00:55.60" lane="1" heatid="5013" />
                <RESULT resultid="598" eventid="10" swimtime="00:00:24.84" lane="1" heatid="10013" />
                <RESULT resultid="599" eventid="12" swimtime="00:01:06.19" lane="8" heatid="12001" />
                <RESULT resultid="600" eventid="13" swimtime="00:02:07.67" lane="5" heatid="13008">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:03.05" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="181" birthdate="2016-01-01" gender="M" lastname="Mund" firstname="Karl" license="0">
              <RESULTS>
                <RESULT resultid="601" eventid="2" swimtime="00:00:41.17" lane="2" heatid="2001" />
                <RESULT resultid="602" eventid="4" status="DSQ" swimtime="00:00:00.00" lane="6" heatid="4001" comment="aufgegeben nach 20 m" />
                <RESULT resultid="603" eventid="7" swimtime="00:00:58.95" lane="3" heatid="7001" />
                <RESULT resultid="604" eventid="11" swimtime="00:00:53.47" lane="8" heatid="11001" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="182" birthdate="2011-01-01" gender="F" lastname="Döll" firstname="Katharina Martha" license="0">
              <RESULTS>
                <RESULT resultid="605" eventid="3" status="DSQ" swimtime="00:06:13.30" lane="3" heatid="3004" comment="Falscher Start.">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:19.41" />
                    <SPLIT distance="200" swimtime="00:02:58.37" />
                    <SPLIT distance="300" swimtime="00:04:37.64" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="606" eventid="5" swimtime="00:01:16.94" lane="5" heatid="5004" />
                <RESULT resultid="607" eventid="10" swimtime="00:00:33.00" lane="8" heatid="10004" />
                <RESULT resultid="608" eventid="13" swimtime="00:02:53.87" lane="7" heatid="13006">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:19.68" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="184" birthdate="2010-01-01" gender="M" lastname="Hochstein" firstname="Maddox Lee" license="0">
              <RESULTS>
                <RESULT resultid="614" eventid="3" swimtime="00:05:00.07" lane="4" heatid="3005">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:08.90" />
                    <SPLIT distance="200" swimtime="00:02:28.44" />
                    <SPLIT distance="300" swimtime="00:03:48.30" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="615" eventid="5" swimtime="00:01:02.39" lane="1" heatid="5011" />
                <RESULT resultid="616" eventid="10" swimtime="00:00:26.88" lane="1" heatid="10011" />
                <RESULT resultid="617" eventid="13" swimtime="00:02:25.20" lane="6" heatid="13008">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:10.09" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="185" birthdate="2009-01-01" gender="F" lastname="Blumenstein" firstname="Martha" license="0">
              <RESULTS>
                <RESULT resultid="618" eventid="1" swimtime="00:00:24.71" lane="8" heatid="1003" />
                <RESULT resultid="619" eventid="3" swimtime="00:04:37.35" lane="5" heatid="3007">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:05.96" />
                    <SPLIT distance="200" swimtime="00:02:18.04" />
                    <SPLIT distance="300" swimtime="00:03:30.63" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="620" eventid="5" swimtime="00:00:54.96" lane="6" heatid="5014" />
                <RESULT resultid="621" eventid="10" swimtime="00:00:25.06" lane="3" heatid="10013" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="186" birthdate="2012-01-01" gender="F" lastname="Palchyk" firstname="Myroslava" license="0">
              <RESULTS>
                <RESULT resultid="622" eventid="5" swimtime="00:01:03.64" lane="1" heatid="5010" />
                <RESULT resultid="623" eventid="8" swimtime="00:00:29.91" lane="3" heatid="8004" />
                <RESULT resultid="624" eventid="10" swimtime="00:00:28.09" lane="5" heatid="10009" />
                <RESULT resultid="625" eventid="13" swimtime="00:02:24.10" lane="3" heatid="13007">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:12.98" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="187" birthdate="2012-01-01" gender="F" lastname="Schulze" firstname="Paula" license="0">
              <RESULTS>
                <RESULT resultid="626" eventid="5" swimtime="00:01:12.04" lane="3" heatid="5006" />
                <RESULT resultid="627" eventid="8" swimtime="00:00:35.73" lane="7" heatid="8004" />
                <RESULT resultid="628" eventid="10" swimtime="00:00:31.92" lane="6" heatid="10005" />
                <RESULT resultid="629" eventid="13" swimtime="00:02:45.60" lane="5" heatid="13005">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:17.78" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY number="1" gender="X" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="559" eventid="14" swimtime="00:02:40.26" lane="1" heatid="14003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:49.35" />
                    <SPLIT distance="200" swimtime="00:01:46.48" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="172" number="1" />
                    <RELAYPOSITION athleteid="179" number="2" />
                    <RELAYPOSITION athleteid="171" number="3" />
                    <RELAYPOSITION athleteid="185" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" gender="X" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="560" eventid="14" swimtime="00:02:54.77" lane="3" heatid="14002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:52.46" />
                    <SPLIT distance="200" swimtime="00:01:52.06" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="173" number="1" />
                    <RELAYPOSITION athleteid="177" number="2" />
                    <RELAYPOSITION athleteid="180" number="3" />
                    <RELAYPOSITION athleteid="187" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" gender="X" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="561" eventid="14" swimtime="00:03:07.47" lane="6" heatid="14001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:58.20" />
                    <SPLIT distance="200" swimtime="00:02:01.56" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="178" number="1" />
                    <RELAYPOSITION athleteid="184" number="2" />
                    <RELAYPOSITION athleteid="186" number="3" />
                    <RELAYPOSITION athleteid="174" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB name="TC Chemie Greiz e.V." nation="GER" region="35" code="174117">
          <ATHLETES>
            <ATHLETE athleteid="58" birthdate="2009-01-01" gender="F" lastname="Naupold" firstname="Celina" license="0">
              <RESULTS>
                <RESULT resultid="193" eventid="1" swimtime="00:00:22.74" lane="6" heatid="1003" />
                <RESULT resultid="194" eventid="5" swimtime="00:00:53.97" lane="6" heatid="5013" />
                <RESULT resultid="195" eventid="10" swimtime="00:00:24.59" lane="2" heatid="10012" />
                <RESULT resultid="196" eventid="12" swimtime="00:00:55.97" lane="3" heatid="12003" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="59" birthdate="2011-01-01" gender="F" lastname="Brendel" firstname="Emma" license="0">
              <RESULTS>
                <RESULT resultid="197" eventid="5" swimtime="00:00:55.58" lane="7" heatid="5013" />
                <RESULT resultid="198" eventid="10" swimtime="00:00:24.66" lane="2" heatid="10013" />
                <RESULT resultid="199" eventid="12" swimtime="00:00:58.87" lane="7" heatid="12003" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="60" birthdate="2011-01-01" gender="F" lastname="Volger" firstname="Eva" license="0">
              <RESULTS>
                <RESULT resultid="200" eventid="3" swimtime="00:05:33.66" lane="8" heatid="3003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:17.47" />
                    <SPLIT distance="200" swimtime="00:02:45.31" />
                    <SPLIT distance="300" swimtime="00:04:12.33" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="201" eventid="5" swimtime="00:01:12.03" lane="3" heatid="5007" />
                <RESULT resultid="202" eventid="10" swimtime="00:00:32.25" lane="2" heatid="10005" />
                <RESULT resultid="203" eventid="13" swimtime="00:02:39.16" lane="4" heatid="13005">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:15.38" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="61" birthdate="2008-01-01" gender="M" lastname="Lose" firstname="Fabian" license="0">
              <RESULTS>
                <RESULT resultid="204" eventid="3" swimtime="00:04:45.28" lane="5" heatid="3006">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:04.46" />
                    <SPLIT distance="200" swimtime="00:02:19.23" />
                    <SPLIT distance="300" swimtime="00:03:36.55" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="205" eventid="5" status="DSQ" swimtime="00:00:00.00" lane="7" heatid="5012" comment="falsche Ausrüstung (Flosse beim Start verloren)&#xA;aufgegeben nach 3 m&#xA;" />
                <RESULT resultid="206" eventid="10" swimtime="00:00:26.35" lane="2" heatid="10011" />
                <RESULT resultid="207" eventid="13" swimtime="00:02:10.58" lane="4" heatid="13008">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:02.77" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="64" birthdate="2008-01-01" gender="M" lastname="Robenz" firstname="Jean Robin" license="0">
              <RESULTS>
                <RESULT resultid="210" eventid="1" status="DSQ" swimtime="00:00:21.23" lane="2" heatid="1003" comment="falscher Start" />
                <RESULT resultid="211" eventid="5" swimtime="00:00:50.91" lane="3" heatid="5013" />
                <RESULT resultid="212" eventid="10" swimtime="00:00:22.45" lane="3" heatid="10015" />
                <RESULT resultid="213" eventid="12" status="DSQ" swimtime="00:00:49.09" lane="1" heatid="12004" comment="Falscher Start.." />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="65" birthdate="2014-01-01" gender="F" lastname="Zeil" firstname="Johanna" license="0">
              <RESULTS>
                <RESULT resultid="214" eventid="5" swimtime="00:01:42.54" lane="6" heatid="5001" />
                <RESULT resultid="215" eventid="8" status="DSQ" swimtime="00:00:49.05" lane="2" heatid="8001" comment="Falscher Schwimmstil. &#xA;Mehrere Wechselbeinschläge nach dem Start." />
                <RESULT resultid="216" eventid="10" swimtime="00:00:43.43" lane="6" heatid="10001" />
                <RESULT resultid="217" eventid="13" swimtime="00:03:46.10" lane="3" heatid="13001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:44.68" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="67" birthdate="2015-01-01" gender="M" lastname="Schulze" firstname="Joshua" license="0">
              <RESULTS>
                <RESULT resultid="221" eventid="2" swimtime="00:00:35.88" lane="3" heatid="2002" />
                <RESULT resultid="222" eventid="4" swimtime="00:00:16.75" lane="3" heatid="4001" />
                <RESULT resultid="643" eventid="5" swimtime="00:01:18.95" lane="6" heatid="5003" />
                <RESULT resultid="223" eventid="7" swimtime="00:00:36.59" lane="3" heatid="7002" />
                <RESULT resultid="644" eventid="10" swimtime="00:00:37.61" lane="6" heatid="10002" />
                <RESULT resultid="650" eventid="11" swimtime="00:00:41.33" lane="3" heatid="11001" />
                <RESULT resultid="645" eventid="13" swimtime="00:02:55.93" lane="7" heatid="13003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:25.01" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="69" birthdate="2009-01-01" gender="M" lastname="Heydel" firstname="Linus" license="0">
              <RESULTS>
                <RESULT resultid="228" eventid="1" swimtime="00:00:20.96" lane="3" heatid="1004" />
                <RESULT resultid="229" eventid="3" swimtime="00:04:13.04" lane="5" heatid="3008">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:56.36" />
                    <SPLIT distance="200" swimtime="00:02:01.86" />
                    <SPLIT distance="300" swimtime="00:03:10.45" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="230" eventid="6" swimtime="00:04:42.08" lane="6" heatid="6001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:01.01" />
                    <SPLIT distance="200" swimtime="00:02:12.82" />
                    <SPLIT distance="300" swimtime="00:03:30.31" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="231" eventid="12" swimtime="00:00:52.42" lane="5" heatid="12003" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="70" birthdate="2011-01-01" gender="F" lastname="Leonhardt" firstname="Ronja" license="0">
              <RESULTS>
                <RESULT resultid="232" eventid="3" swimtime="00:05:18.10" lane="2" heatid="3005">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:13.45" />
                    <SPLIT distance="200" swimtime="00:02:38.15" />
                    <SPLIT distance="300" swimtime="00:04:01.43" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="233" eventid="5" swimtime="00:01:09.13" lane="8" heatid="5009" />
                <RESULT resultid="234" eventid="10" swimtime="00:00:31.44" lane="2" heatid="10007" />
                <RESULT resultid="235" eventid="13" swimtime="00:02:31.45" lane="4" heatid="13007">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:14.51" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="71" birthdate="2011-01-01" gender="F" lastname="Klar" firstname="Sophia" license="0">
              <RESULTS>
                <RESULT resultid="236" eventid="3" swimtime="00:06:22.67" lane="3" heatid="3001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:25.82" />
                    <SPLIT distance="200" swimtime="00:03:09.98" />
                    <SPLIT distance="300" swimtime="00:04:47.52" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="237" eventid="5" swimtime="00:01:12.62" lane="1" heatid="5007" />
                <RESULT resultid="238" eventid="10" swimtime="00:00:30.12" lane="7" heatid="10008" />
                <RESULT resultid="239" eventid="12" swimtime="00:01:13.72" lane="2" heatid="12001" />
                <RESULT resultid="240" eventid="13" swimtime="00:03:04.76" lane="2" heatid="13003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:31.97" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="73" birthdate="2016-01-01" gender="M" lastname="Hierold" firstname="Theodor" license="0">
              <RESULTS>
                <RESULT resultid="243" eventid="2" swimtime="00:00:38.47" lane="2" heatid="2002" />
                <RESULT resultid="641" eventid="5" swimtime="00:01:25.80" lane="7" heatid="5002" />
                <RESULT resultid="244" eventid="7" swimtime="00:00:39.20" lane="6" heatid="7002" />
                <RESULT resultid="642" eventid="10" swimtime="00:00:39.75" lane="1" heatid="10002" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="74" birthdate="2014-01-01" gender="M" lastname="Volger" firstname="Tom" license="0">
              <RESULTS>
                <RESULT resultid="245" eventid="3" swimtime="00:05:44.35" lane="4" heatid="3002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:19.97" />
                    <SPLIT distance="200" swimtime="00:02:48.02" />
                    <SPLIT distance="300" swimtime="00:04:18.44" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="246" eventid="5" swimtime="00:01:15.18" lane="2" heatid="5005" />
                <RESULT resultid="247" eventid="8" swimtime="00:00:37.58" lane="5" heatid="8003" />
                <RESULT resultid="248" eventid="10" swimtime="00:00:34.48" lane="7" heatid="10004" />
                <RESULT resultid="249" eventid="13" swimtime="00:02:46.34" lane="8" heatid="13006">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:19.72" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="75" birthdate="2012-01-01" gender="M" lastname="Sochynskyi" firstname="Vadym" license="0">
              <RESULTS>
                <RESULT resultid="250" eventid="3" swimtime="00:05:16.01" lane="7" heatid="3005">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:12.78" />
                    <SPLIT distance="200" swimtime="00:02:34.05" />
                    <SPLIT distance="300" swimtime="00:03:57.77" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="251" eventid="5" swimtime="00:01:05.67" lane="3" heatid="5009" />
                <RESULT resultid="252" eventid="8" swimtime="00:00:31.22" lane="6" heatid="8004" />
                <RESULT resultid="253" eventid="10" swimtime="00:00:29.14" lane="2" heatid="10008" />
                <RESULT resultid="254" eventid="12" swimtime="00:01:19.32" lane="1" heatid="12002" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="76" birthdate="2016-01-01" gender="F" lastname="Volger" firstname="Lea" license="0">
              <RESULTS>
                <RESULT resultid="255" eventid="5" status="DSQ" swimtime="00:01:22.41" lane="8" heatid="5003" comment="Falscher Start" />
                <RESULT resultid="256" eventid="10" swimtime="00:00:36.74" lane="5" heatid="10002" />
                <RESULT resultid="257" eventid="13" swimtime="00:03:02.53" lane="5" heatid="13002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:26.22" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY number="1" gender="X" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="208" eventid="14" swimtime="00:02:39.16" lane="8" heatid="14003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:49.33" />
                    <SPLIT distance="200" swimtime="00:01:45.08" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="64" number="1" />
                    <RELAYPOSITION athleteid="59" number="2" />
                    <RELAYPOSITION athleteid="58" number="3" />
                    <RELAYPOSITION athleteid="61" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" gender="X" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="209" eventid="14" swimtime="00:03:11.51" lane="8" heatid="14002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:55.05" />
                    <SPLIT distance="200" swimtime="00:02:04.68" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="69" number="1" />
                    <RELAYPOSITION athleteid="70" number="2" />
                    <RELAYPOSITION athleteid="75" number="3" />
                    <RELAYPOSITION athleteid="60" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB name="TC fez Berlin" nation="GER" region="21" code="0">
          <ATHLETES>
            <ATHLETE athleteid="119" birthdate="2014-01-01" gender="M" lastname="Bowe" firstname="Constantin" license="0">
              <RESULTS>
                <RESULT resultid="369" eventid="5" swimtime="00:01:18.05" lane="5" heatid="5002" />
                <RESULT resultid="370" eventid="8" swimtime="00:00:38.31" lane="6" heatid="8003" />
                <RESULT resultid="371" eventid="10" swimtime="00:00:34.83" lane="3" heatid="10002" />
                <RESULT resultid="372" eventid="13" swimtime="00:03:03.35" lane="4" heatid="13002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:28.70" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="120" birthdate="2015-01-01" gender="F" lastname="Just" firstname="Elsa" license="0">
              <RESULTS>
                <RESULT resultid="373" eventid="2" swimtime="00:00:40.75" lane="1" heatid="2002" />
                <RESULT resultid="374" eventid="4" status="DSQ" swimtime="00:00:00.00" lane="5" heatid="4001" comment="aufgegeben nach 20 m" />
                <RESULT resultid="638" eventid="5" swimtime="00:01:33.75" lane="2" heatid="5002" />
                <RESULT resultid="375" eventid="7" swimtime="00:00:44.97" lane="5" heatid="7002" />
                <RESULT resultid="376" eventid="11" swimtime="00:00:43.95" lane="4" heatid="11001" />
                <RESULT resultid="639" eventid="13" swimtime="00:03:11.92" lane="4" heatid="13001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:32.96" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="121" birthdate="2006-01-01" gender="M" lastname="Schlobohm" firstname="Enrico" license="0">
              <RESULTS>
                <RESULT resultid="377" eventid="1" swimtime="00:00:17.78" lane="2" heatid="1007" />
                <RESULT resultid="378" eventid="5" swimtime="00:00:42.53" lane="5" heatid="5018" />
                <RESULT resultid="379" eventid="10" swimtime="00:00:19.58" lane="2" heatid="10018" />
                <RESULT resultid="380" eventid="12" swimtime="00:00:45.27" lane="7" heatid="12005" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="122" birthdate="2005-01-01" gender="F" lastname="Tesch" firstname="Florentine" license="0">
              <RESULTS>
                <RESULT resultid="381" eventid="1" swimtime="00:00:18.75" lane="8" heatid="1007" />
                <RESULT resultid="382" eventid="5" swimtime="00:00:46.27" lane="5" heatid="5017" />
                <RESULT resultid="383" eventid="6" status="DSQ" swimtime="00:00:00.00" lane="5" heatid="6001" comment="Gesicht aus dem Wasser bei 190 m.">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:57.02" />
                    <SPLIT distance="200" swimtime="00:02:17.52" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="384" eventid="10" swimtime="00:00:19.66" lane="6" heatid="10017" />
                <RESULT resultid="385" eventid="12" swimtime="00:00:45.96" lane="7" heatid="12004" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="123" birthdate="2014-01-01" gender="F" lastname="Rüdiger" firstname="Henrikje" license="0">
              <RESULTS>
                <RESULT resultid="386" eventid="3" swimtime="00:06:32.34" lane="8" heatid="3002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:29.68" />
                    <SPLIT distance="200" swimtime="00:03:12.91" />
                    <SPLIT distance="300" swimtime="00:05:00.95" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="387" eventid="5" swimtime="00:01:16.51" lane="7" heatid="5006" />
                <RESULT resultid="388" eventid="8" swimtime="00:00:38.81" lane="2" heatid="8003" />
                <RESULT resultid="389" eventid="10" swimtime="00:00:33.46" lane="1" heatid="10004" />
                <RESULT resultid="390" eventid="13" swimtime="00:02:55.70" lane="3" heatid="13004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:26.17" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="124" birthdate="2011-01-01" gender="M" lastname="Bardo" firstname="John" license="0">
              <RESULTS>
                <RESULT resultid="391" eventid="5" swimtime="00:01:23.01" lane="2" heatid="5003" />
                <RESULT resultid="392" eventid="10" swimtime="00:00:34.97" lane="2" heatid="10003" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="125" birthdate="2013-01-01" gender="F" lastname="Harder" firstname="Juli" license="0">
              <RESULTS>
                <RESULT resultid="393" eventid="3" swimtime="00:05:55.27" lane="7" heatid="3002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:24.32" />
                    <SPLIT distance="200" swimtime="00:02:55.88" />
                    <SPLIT distance="300" swimtime="00:04:29.78" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="394" eventid="5" swimtime="00:01:27.95" lane="6" heatid="5004" />
                <RESULT resultid="395" eventid="8" swimtime="00:00:40.58" lane="3" heatid="8003" />
                <RESULT resultid="396" eventid="10" swimtime="00:00:36.94" lane="1" heatid="10003" />
                <RESULT resultid="397" eventid="13" swimtime="00:03:02.72" lane="7" heatid="13005">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:31.17" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="127" birthdate="2007-01-01" gender="F" lastname="Schikora" firstname="Luise" license="0">
              <RESULTS>
                <RESULT resultid="403" eventid="1" swimtime="00:00:20.04" lane="7" heatid="1006" />
                <RESULT resultid="404" eventid="5" swimtime="00:00:48.83" lane="7" heatid="5017" />
                <RESULT resultid="405" eventid="10" status="DNS" swimtime="00:00:00.00" lane="6" heatid="10016" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="128" birthdate="2007-01-01" gender="F" lastname="Rüdiger" firstname="Marielena" license="0">
              <RESULTS>
                <RESULT resultid="406" eventid="3" swimtime="00:04:41.92" lane="3" heatid="3006">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:09.54" />
                    <SPLIT distance="200" swimtime="00:02:25.18" />
                    <SPLIT distance="300" swimtime="00:03:36.13" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="407" eventid="5" status="DSQ" swimtime="00:00:57.74" lane="4" heatid="5012" comment="Tauchzüge außerhalb der 15m-Zonen (mehrere Tauchzüge außerhalb der 15m-Zone)" />
                <RESULT resultid="408" eventid="10" swimtime="00:00:26.04" lane="6" heatid="10011" />
                <RESULT resultid="409" eventid="12" swimtime="00:00:58.54" lane="8" heatid="12003" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="129" birthdate="2013-01-01" gender="F" lastname="Volkert" firstname="Sophia" license="0">
              <RESULTS>
                <RESULT resultid="410" eventid="5" swimtime="00:01:18.69" lane="5" heatid="5003" />
                <RESULT resultid="411" eventid="8" swimtime="00:00:39.39" lane="7" heatid="8003" />
                <RESULT resultid="412" eventid="10" swimtime="00:00:34.94" lane="7" heatid="10003" />
                <RESULT resultid="413" eventid="13" swimtime="00:03:02.17" lane="3" heatid="13003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:27.69" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="130" birthdate="2013-01-01" gender="F" lastname="Ringling" firstname="Sophie" license="0">
              <RESULTS>
                <RESULT resultid="414" eventid="3" swimtime="00:05:36.04" lane="6" heatid="3003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:19.46" />
                    <SPLIT distance="200" swimtime="00:02:46.47" />
                    <SPLIT distance="300" swimtime="00:04:14.02" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="415" eventid="5" swimtime="00:01:16.12" lane="6" heatid="5005" />
                <RESULT resultid="416" eventid="8" swimtime="00:00:36.34" lane="8" heatid="8004" />
                <RESULT resultid="417" eventid="10" swimtime="00:00:33.88" lane="7" heatid="10005" />
                <RESULT resultid="418" eventid="13" swimtime="00:02:52.22" lane="6" heatid="13005">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:23.58" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="191" birthdate="2012-01-01" gender="F" lastname="Lukaschewska" firstname="Elena" license="0">
              <RESULTS>
                <RESULT resultid="646" eventid="3" status="DSQ" swimtime="00:05:57.02" lane="8" heatid="3004" comment="Falsche Ausrüstung (Flosse verloren bei 200m)">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:15.55" />
                    <SPLIT distance="200" swimtime="00:02:46.23" />
                    <SPLIT distance="300" swimtime="00:04:29.62" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="647" eventid="5" swimtime="00:01:16.88" lane="4" heatid="5004" />
                <RESULT resultid="648" eventid="10" status="DSQ" swimtime="00:00:33.23" lane="5" heatid="10007" comment="falscher Start" />
                <RESULT resultid="649" eventid="13" swimtime="00:02:52.19" lane="5" heatid="13004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:21.41" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY number="1" gender="X" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="366" eventid="14" swimtime="00:03:11.64" lane="7" heatid="14003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:56.20" />
                    <SPLIT distance="200" swimtime="00:02:04.63" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="122" number="1" />
                    <RELAYPOSITION athleteid="191" number="2" />
                    <RELAYPOSITION athleteid="128" number="3" />
                    <RELAYPOSITION athleteid="129" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="2" gender="X" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="367" eventid="14" swimtime="00:03:46.85" lane="4" heatid="14001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:55.73" />
                    <SPLIT distance="200" swimtime="00:02:22.06" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="121" number="1" />
                    <RELAYPOSITION athleteid="130" number="2" />
                    <RELAYPOSITION athleteid="123" number="3" />
                    <RELAYPOSITION athleteid="120" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="3" gender="X" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="368" eventid="14" swimtime="00:03:42.01" lane="3" heatid="14001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:57.51" />
                    <SPLIT distance="200" swimtime="00:02:21.06" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="127" number="1" />
                    <RELAYPOSITION athleteid="125" number="2" />
                    <RELAYPOSITION athleteid="119" number="3" />
                    <RELAYPOSITION athleteid="124" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB name="TC Harz" nation="GER" region="27" code="0">
          <ATHLETES>
            <ATHLETE athleteid="137" birthdate="2011-01-01" gender="M" lastname="Beier" firstname="Anton" license="0">
              <RESULTS>
                <RESULT resultid="433" eventid="3" swimtime="00:04:51.07" lane="7" heatid="3006">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:11.47" />
                    <SPLIT distance="200" swimtime="00:02:27.14" />
                    <SPLIT distance="300" swimtime="00:03:41.10" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="434" eventid="5" status="DSQ" swimtime="00:01:05.03" lane="3" heatid="5010" comment="falscher Start" />
                <RESULT resultid="435" eventid="10" status="DSQ" swimtime="00:00:29.08" lane="1" heatid="10010" comment="Tauchzüger außerhalb der 15m-Zone bei ca 20 m" />
                <RESULT resultid="436" eventid="13" swimtime="00:02:21.52" lane="8" heatid="13008">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:10.24" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="138" birthdate="2014-01-01" gender="M" lastname="Hass" firstname="Ben Henry" license="0">
              <RESULTS>
                <RESULT resultid="437" eventid="3" swimtime="00:05:39.66" lane="1" heatid="3004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:21.35" />
                    <SPLIT distance="200" swimtime="00:02:49.59" />
                    <SPLIT distance="300" swimtime="00:04:19.98" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="438" eventid="5" swimtime="00:01:23.30" lane="8" heatid="5008" />
                <RESULT resultid="439" eventid="10" swimtime="00:00:32.89" lane="1" heatid="10007" />
                <RESULT resultid="440" eventid="13" swimtime="00:02:43.15" lane="7" heatid="13007">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:20.93" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="139" birthdate="2007-01-01" gender="F" lastname="Risse" firstname="Elisabeth" license="0">
              <RESULTS>
                <RESULT resultid="441" eventid="1" swimtime="00:00:22.32" lane="6" heatid="1004" />
                <RESULT resultid="442" eventid="3" swimtime="00:04:26.48" lane="7" heatid="3009">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:01.27" />
                    <SPLIT distance="200" swimtime="00:02:09.31" />
                    <SPLIT distance="300" swimtime="00:03:18.76" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="443" eventid="5" swimtime="00:00:54.49" lane="1" heatid="5016" />
                <RESULT resultid="444" eventid="10" swimtime="00:00:23.48" lane="8" heatid="10016" />
                <RESULT resultid="445" eventid="13" swimtime="00:02:03.37" lane="5" heatid="13011">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:57.88" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="140" birthdate="2012-01-01" gender="M" lastname="Rolle" firstname="Emilius" license="0">
              <RESULTS>
                <RESULT resultid="446" eventid="3" swimtime="00:05:39.88" lane="1" heatid="3002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:17.06" />
                    <SPLIT distance="200" swimtime="00:02:47.46" />
                    <SPLIT distance="300" swimtime="00:04:16.96" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="447" eventid="5" swimtime="00:01:10.43" lane="7" heatid="5008" />
                <RESULT resultid="448" eventid="10" swimtime="00:00:28.78" lane="1" heatid="10008" />
                <RESULT resultid="449" eventid="13" swimtime="00:02:41.79" lane="6" heatid="13003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:17.96" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="141" birthdate="2011-01-01" gender="F" lastname="Chyla" firstname="Emma" license="0">
              <RESULTS>
                <RESULT resultid="450" eventid="3" status="DSQ" swimtime="00:06:05.86" lane="3" heatid="3002" comment="Falscher Start.">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:24.75" />
                    <SPLIT distance="200" swimtime="00:03:01.95" />
                    <SPLIT distance="300" swimtime="00:04:38.43" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="451" eventid="5" swimtime="00:01:11.89" lane="5" heatid="5007" />
                <RESULT resultid="452" eventid="10" swimtime="00:00:30.82" lane="3" heatid="10006" />
                <RESULT resultid="453" eventid="13" status="DSQ" swimtime="00:02:46.80" lane="8" heatid="13005" comment="Tauchzüge außerhalb der 15m-Zonen bei ca 125 m">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:17.72" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="142" birthdate="2012-01-01" gender="M" lastname="Neumann" firstname="Erik" license="0">
              <RESULTS>
                <RESULT resultid="454" eventid="3" swimtime="00:05:20.22" lane="2" heatid="3004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:13.52" />
                    <SPLIT distance="200" swimtime="00:02:36.49" />
                    <SPLIT distance="300" swimtime="00:04:01.24" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="455" eventid="5" swimtime="00:01:08.68" lane="6" heatid="5008" />
                <RESULT resultid="456" eventid="10" swimtime="00:00:31.68" lane="6" heatid="10006" />
                <RESULT resultid="457" eventid="13" swimtime="00:02:34.79" lane="2" heatid="13006">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:16.85" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="143" birthdate="2014-01-01" gender="F" lastname="Brüser" firstname="Fina Maria" license="0">
              <RESULTS>
                <RESULT resultid="458" eventid="5" swimtime="00:01:24.93" lane="6" heatid="5002" />
                <RESULT resultid="459" eventid="8" swimtime="00:00:41.23" lane="4" heatid="8002" />
                <RESULT resultid="460" eventid="10" swimtime="00:00:38.84" lane="6" heatid="10003" />
                <RESULT resultid="461" eventid="13" swimtime="00:03:08.77" lane="6" heatid="13002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:30.03" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="144" birthdate="2014-01-01" gender="M" lastname="Klinner" firstname="Floris" license="0">
              <RESULTS>
                <RESULT resultid="462" eventid="5" swimtime="00:01:22.56" lane="7" heatid="5004" />
                <RESULT resultid="463" eventid="8" swimtime="00:00:37.47" lane="5" heatid="8002" />
                <RESULT resultid="464" eventid="10" swimtime="00:00:37.03" lane="5" heatid="10003" />
                <RESULT resultid="465" eventid="13" swimtime="00:03:06.34" lane="8" heatid="13003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:31.20" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="145" birthdate="2012-01-01" gender="F" lastname="Dieck" firstname="Franziska" license="0">
              <RESULTS>
                <RESULT resultid="466" eventid="3" status="DSQ" swimtime="00:05:51.80" lane="5" heatid="3002" comment="Falscher Start,">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:19.82" />
                    <SPLIT distance="200" swimtime="00:02:50.94" />
                    <SPLIT distance="300" swimtime="00:04:22.34" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="467" eventid="5" swimtime="00:01:17.23" lane="4" heatid="5005" />
                <RESULT resultid="468" eventid="10" swimtime="00:00:31.39" lane="5" heatid="10005" />
                <RESULT resultid="469" eventid="13" swimtime="00:02:50.10" lane="6" heatid="13004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:20.85" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="146" birthdate="2008-01-01" gender="M" lastname="Härter" firstname="Fynn" license="0">
              <RESULTS>
                <RESULT resultid="470" eventid="1" swimtime="00:00:20.04" lane="7" heatid="1005" />
                <RESULT resultid="471" eventid="3" swimtime="00:03:59.25" lane="6" heatid="3009">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:54.77" />
                    <SPLIT distance="200" swimtime="00:01:56.89" />
                    <SPLIT distance="300" swimtime="00:03:00.58" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="472" eventid="5" swimtime="00:00:50.31" lane="8" heatid="5016" />
                <RESULT resultid="473" eventid="10" swimtime="00:00:27.09" lane="7" heatid="10016" />
                <RESULT resultid="474" eventid="13" swimtime="00:01:52.57" lane="1" heatid="13012">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:52.75" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="147" birthdate="2011-01-01" gender="F" lastname="Dachner" firstname="Helena" license="0">
              <RESULTS>
                <RESULT resultid="475" eventid="3" status="DNS" swimtime="00:00:00.00" lane="2" heatid="3003" />
                <RESULT resultid="476" eventid="5" status="DNS" swimtime="00:00:00.00" lane="1" heatid="5004" />
                <RESULT resultid="477" eventid="10" status="DNS" swimtime="00:00:00.00" lane="4" heatid="10004" />
                <RESULT resultid="478" eventid="13" status="DNS" swimtime="00:00:00.00" lane="5" heatid="13003" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="148" birthdate="2011-01-01" gender="F" lastname="Langer" firstname="Ida" license="0">
              <RESULTS>
                <RESULT resultid="479" eventid="3" swimtime="00:05:37.53" lane="3" heatid="3003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:18.33" />
                    <SPLIT distance="200" swimtime="00:02:46.45" />
                    <SPLIT distance="300" swimtime="00:04:14.36" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="480" eventid="5" swimtime="00:01:25.10" lane="4" heatid="5007" />
                <RESULT resultid="481" eventid="10" swimtime="00:00:31.68" lane="7" heatid="10006" />
                <RESULT resultid="482" eventid="13" swimtime="00:02:37.78" lane="8" heatid="13004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:12.71" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="149" birthdate="2004-01-01" gender="M" lastname="Hass" firstname="Jan Henrik" license="0">
              <RESULTS>
                <RESULT resultid="483" eventid="1" swimtime="00:00:17.59" lane="7" heatid="1007" />
                <RESULT resultid="484" eventid="5" swimtime="00:00:43.50" lane="2" heatid="5018" />
                <RESULT resultid="485" eventid="10" swimtime="00:00:19.63" lane="3" heatid="10018" />
                <RESULT resultid="486" eventid="13" swimtime="00:01:43.90" lane="3" heatid="13012">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:49.00" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="150" birthdate="2012-01-01" gender="F" lastname="Krzizak" firstname="Lana" license="0">
              <RESULTS>
                <RESULT resultid="487" eventid="3" swimtime="00:05:55.99" lane="4" heatid="3001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:21.35" />
                    <SPLIT distance="200" swimtime="00:02:55.55" />
                    <SPLIT distance="300" swimtime="00:04:30.05" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="488" eventid="5" swimtime="00:01:15.38" lane="8" heatid="5007" />
                <RESULT resultid="489" eventid="10" swimtime="00:00:32.28" lane="4" heatid="10005" />
                <RESULT resultid="490" eventid="13" swimtime="00:02:56.69" lane="2" heatid="13005">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:25.39" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="151" birthdate="2003-01-01" gender="M" lastname="von Gynz Rekowski" firstname="Louis" license="0">
              <RESULTS>
                <RESULT resultid="491" eventid="1" status="DSQ" swimtime="00:00:20.67" lane="6" heatid="1005" comment="falscher Start" />
                <RESULT resultid="492" eventid="5" swimtime="00:00:55.72" lane="3" heatid="5016" />
                <RESULT resultid="493" eventid="10" status="DSQ" swimtime="00:00:25.00" lane="4" heatid="10016" comment="Tauchzüge außerhalb der 15m-Zone bei ca. 20 m" />
                <RESULT resultid="494" eventid="12" swimtime="00:00:51.81" lane="1" heatid="12005" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="152" birthdate="2009-01-01" gender="F" lastname="Zündel" firstname="Marlene" license="0">
              <RESULTS>
                <RESULT resultid="495" eventid="1" swimtime="00:00:22.16" lane="7" heatid="1003" />
                <RESULT resultid="496" eventid="3" swimtime="00:04:31.05" lane="2" heatid="3008">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:02.61" />
                    <SPLIT distance="200" swimtime="00:02:14.37" />
                    <SPLIT distance="300" swimtime="00:03:24.37" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="497" eventid="5" swimtime="00:00:55.09" lane="8" heatid="5015" />
                <RESULT resultid="498" eventid="10" swimtime="00:00:24.00" lane="3" heatid="10014" />
                <RESULT resultid="499" eventid="13" status="DSQ" swimtime="00:02:01.73" lane="8" heatid="13011" comment="Falscher Start.&#xA;Tauchzüge außerhalb der 15m-Zonen bei ca. 40 m.">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:56.31" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="153" birthdate="2008-01-01" gender="F" lastname="Weißenborn" firstname="Marnie" license="0">
              <RESULTS>
                <RESULT resultid="500" eventid="1" swimtime="00:00:20.50" lane="5" heatid="1005" />
                <RESULT resultid="501" eventid="3" swimtime="00:04:07.53" lane="3" heatid="3009">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:56.69" />
                    <SPLIT distance="200" swimtime="00:02:00.19" />
                    <SPLIT distance="300" swimtime="00:03:04.75" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="502" eventid="5" swimtime="00:00:48.91" lane="2" heatid="5017" />
                <RESULT resultid="503" eventid="10" swimtime="00:00:22.14" lane="3" heatid="10016" />
                <RESULT resultid="504" eventid="13" swimtime="00:01:50.53" lane="6" heatid="13012">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:52.84" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="154" birthdate="2009-01-01" gender="M" lastname="Schmidt" firstname="Matty" license="0">
              <RESULTS>
                <RESULT resultid="505" eventid="1" status="DSQ" swimtime="00:00:00.00" lane="8" heatid="1002" comment="Aufgabe nach 0 m" />
                <RESULT resultid="506" eventid="3" swimtime="00:04:22.57" lane="7" heatid="3008">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:02.20" />
                    <SPLIT distance="200" swimtime="00:02:11.69" />
                    <SPLIT distance="300" swimtime="00:03:18.38" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="507" eventid="5" swimtime="00:00:56.92" lane="4" heatid="5013" />
                <RESULT resultid="508" eventid="10" swimtime="00:00:26.35" lane="7" heatid="10013" />
                <RESULT resultid="509" eventid="13" swimtime="00:02:03.59" lane="7" heatid="13010">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:02.36" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="155" birthdate="2012-01-01" gender="F" lastname="Wegemer" firstname="Mette" license="0">
              <RESULTS>
                <RESULT resultid="510" eventid="3" swimtime="00:06:37.34" lane="2" heatid="3002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:26.24" />
                    <SPLIT distance="200" swimtime="00:03:10.14" />
                    <SPLIT distance="300" swimtime="00:04:54.59" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="511" eventid="5" swimtime="00:01:22.98" lane="3" heatid="5003" />
                <RESULT resultid="512" eventid="10" status="DSQ" swimtime="00:00:34.15" lane="3" heatid="10004" comment="falscher Start" />
                <RESULT resultid="513" eventid="13" swimtime="00:03:03.51" lane="2" heatid="13004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:25.64" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="156" birthdate="2003-01-01" gender="M" lastname="Dalichow" firstname="Noah" license="0">
              <RESULTS>
                <RESULT resultid="514" eventid="1" swimtime="00:00:17.09" lane="3" heatid="1007" />
                <RESULT resultid="515" eventid="5" status="DSQ" swimtime="00:00:48.61" lane="7" heatid="5018" comment="Tauchzüge außerhalb der 15m-Zonen bei ca 90 Meter" />
                <RESULT resultid="516" eventid="10" swimtime="00:00:19.86" lane="5" heatid="10018" />
                <RESULT resultid="517" eventid="12" swimtime="00:00:40.54" lane="5" heatid="12005" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="158" birthdate="2013-01-01" gender="M" lastname="Hoffmeister" firstname="Oskar" license="0">
              <RESULTS>
                <RESULT resultid="519" eventid="3" swimtime="00:05:12.92" lane="1" heatid="3006">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:12.46" />
                    <SPLIT distance="200" swimtime="00:02:33.16" />
                    <SPLIT distance="300" swimtime="00:03:56.27" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="520" eventid="5" swimtime="00:01:06.73" lane="8" heatid="5010" />
                <RESULT resultid="521" eventid="10" swimtime="00:00:30.08" lane="2" heatid="10009" />
                <RESULT resultid="522" eventid="13" swimtime="00:02:26.89" lane="1" heatid="13008">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:10.84" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="159" birthdate="2015-01-01" gender="F" lastname="Meyer" firstname="Ronja" license="0">
              <RESULTS>
                <RESULT resultid="523" eventid="2" swimtime="00:00:38.23" lane="4" heatid="2002" />
                <RESULT resultid="524" eventid="4" swimtime="00:00:17.85" lane="4" heatid="4001" />
                <RESULT resultid="525" eventid="7" swimtime="00:00:37.03" lane="4" heatid="7002" />
                <RESULT resultid="526" eventid="11" swimtime="00:00:37.39" lane="5" heatid="11001" />
                <RESULT resultid="640" eventid="13" status="DSQ" swimtime="00:03:32.26" lane="3" heatid="13002" comment="Falsche Ausrüstung.&#xA;Flosse beim Start verloren." />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="160" birthdate="2007-01-01" gender="F" lastname="von Gynz Rekowski" firstname="Sophie" license="0">
              <RESULTS>
                <RESULT resultid="527" eventid="1" swimtime="00:00:21.43" lane="2" heatid="1004" />
                <RESULT resultid="528" eventid="3" status="DSQ" swimtime="00:04:41.41" lane="8" heatid="3008" comment="Tauchzüge außerhalb der 15 m-Zonen bei ca. 190 m">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:02.89" />
                    <SPLIT distance="200" swimtime="00:02:12.33" />
                    <SPLIT distance="300" swimtime="00:03:28.55" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="529" eventid="5" swimtime="00:00:54.03" lane="3" heatid="5014" />
                <RESULT resultid="530" eventid="10" swimtime="00:00:24.15" lane="1" heatid="10014" />
                <RESULT resultid="531" eventid="13" status="DSQ" swimtime="00:02:04.58" lane="6" heatid="13010" comment="Tauchzüge außerhalb der 15m- Zonen bei ca. 30 Meter.">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:00.49" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="161" birthdate="2009-01-01" gender="M" lastname="Piorun" firstname="Tariq" license="0">
              <RESULTS>
                <RESULT resultid="532" eventid="3" swimtime="00:05:06.12" lane="1" heatid="3003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:07.51" />
                    <SPLIT distance="200" swimtime="00:02:29.29" />
                    <SPLIT distance="300" swimtime="00:03:50.83" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="533" eventid="5" swimtime="00:01:00.79" lane="7" heatid="5009" />
                <RESULT resultid="534" eventid="10" swimtime="00:00:27.26" lane="8" heatid="10009" />
                <RESULT resultid="535" eventid="13" swimtime="00:02:20.65" lane="1" heatid="13007">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:04.30" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="190" birthdate="2003-01-01" gender="M" lastname="Gerlach" firstname="Ruben" license="0" />
          </ATHLETES>
          <RELAYS>
            <RELAY number="1" gender="X" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="518" eventid="14" status="EXH" swimtime="00:02:09.89" lane="4" heatid="14003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:39.13" />
                    <SPLIT distance="200" swimtime="00:01:23.32" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="156" number="1" />
                    <RELAYPOSITION athleteid="149" number="2" />
                    <RELAYPOSITION athleteid="190" number="3" />
                    <RELAYPOSITION athleteid="151" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" gender="X" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="536" eventid="14" swimtime="00:02:27.47" lane="6" heatid="14003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:47.53" />
                    <SPLIT distance="200" swimtime="00:01:36.89" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="146" number="1" />
                    <RELAYPOSITION athleteid="152" number="2" />
                    <RELAYPOSITION athleteid="153" number="3" />
                    <RELAYPOSITION athleteid="154" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB name="TC Marzahn e.V." nation="GER" region="21" code="0">
          <ATHLETES>
            <ATHLETE athleteid="10" birthdate="2010-01-01" gender="F" lastname="Liedloff" firstname="Amelie" license="0">
              <RESULTS>
                <RESULT resultid="22" eventid="3" swimtime="00:04:19.61" lane="1" heatid="3008">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:00.30" />
                    <SPLIT distance="200" swimtime="00:02:07.34" />
                    <SPLIT distance="300" swimtime="00:03:15.62" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="23" eventid="5" swimtime="00:00:54.80" lane="5" heatid="5014" />
                <RESULT resultid="24" eventid="10" swimtime="00:00:24.59" lane="2" heatid="10014" />
                <RESULT resultid="25" eventid="13" swimtime="00:01:59.77" lane="4" heatid="13010">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:57.33" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="11" birthdate="1965-01-01" gender="M" lastname="Ritzer" firstname="Andre" license="0">
              <RESULTS>
                <RESULT resultid="26" eventid="1" swimtime="00:00:24.00" lane="5" heatid="1002" />
                <RESULT resultid="27" eventid="5" swimtime="00:00:59.38" lane="8" heatid="5011" />
                <RESULT resultid="28" eventid="10" swimtime="00:00:26.62" lane="6" heatid="10010" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="12" birthdate="2010-01-01" gender="M" lastname="Kessel" firstname="Benjamin" license="0">
              <RESULTS>
                <RESULT resultid="29" eventid="5" swimtime="00:01:08.56" lane="5" heatid="5006" />
                <RESULT resultid="30" eventid="10" swimtime="00:00:30.14" lane="1" heatid="10005" />
                <RESULT resultid="31" eventid="13" swimtime="00:02:34.85" lane="6" heatid="13006">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:14.59" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="13" birthdate="2008-01-01" gender="F" lastname="Demmrich" firstname="Ella" license="0">
              <RESULTS>
                <RESULT resultid="32" eventid="1" status="DNS" swimtime="00:00:00.00" lane="7" heatid="1002" />
                <RESULT resultid="33" eventid="3" swimtime="00:04:38.84" lane="2" heatid="3007">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:05.13" />
                    <SPLIT distance="200" swimtime="00:02:18.13" />
                    <SPLIT distance="300" swimtime="00:03:30.47" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="34" eventid="5" swimtime="00:00:56.78" lane="6" heatid="5012" />
                <RESULT resultid="35" eventid="10" swimtime="00:00:25.64" lane="7" heatid="10011" />
                <RESULT resultid="36" eventid="13" swimtime="00:02:04.71" lane="8" heatid="13010">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:58.70" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="14" birthdate="2009-01-01" gender="M" lastname="Kupke" firstname="Emil" license="0">
              <RESULTS>
                <RESULT resultid="37" eventid="1" swimtime="00:00:24.32" lane="4" heatid="1002" />
                <RESULT resultid="38" eventid="5" swimtime="00:00:55.26" lane="2" heatid="5013" />
                <RESULT resultid="39" eventid="10" swimtime="00:00:24.40" lane="8" heatid="10013" />
                <RESULT resultid="40" eventid="13" swimtime="00:02:06.77" lane="2" heatid="13009">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:01.20" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="15" birthdate="2004-01-01" gender="F" lastname="May" firstname="Emilie" license="0">
              <RESULTS>
                <RESULT resultid="41" eventid="1" swimtime="00:00:20.42" lane="2" heatid="1005" />
                <RESULT resultid="42" eventid="5" status="DNS" swimtime="00:00:00.00" lane="8" heatid="5017" />
                <RESULT resultid="43" eventid="6" swimtime="00:03:42.19" lane="4" heatid="6001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:49.12" />
                    <SPLIT distance="200" swimtime="00:01:45.78" />
                    <SPLIT distance="300" swimtime="00:02:44.76" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="44" eventid="12" swimtime="00:00:45.43" lane="4" heatid="12004" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="16" birthdate="2009-01-01" gender="M" lastname="Müller" firstname="Erik" license="0">
              <RESULTS>
                <RESULT resultid="45" eventid="5" swimtime="00:01:02.61" lane="2" heatid="5011" />
                <RESULT resultid="46" eventid="10" swimtime="00:00:25.87" lane="3" heatid="10011" />
                <RESULT resultid="47" eventid="13" swimtime="00:02:24.37" lane="3" heatid="13008">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:08.22" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="17" birthdate="2005-01-01" gender="F" lastname="Newerla" firstname="Felicia" license="0">
              <RESULTS>
                <RESULT resultid="48" eventid="1" swimtime="00:00:20.81" lane="1" heatid="1004" />
                <RESULT resultid="49" eventid="5" swimtime="00:00:50.20" lane="1" heatid="5015" />
                <RESULT resultid="50" eventid="10" swimtime="00:00:22.61" lane="5" heatid="10014" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="18" birthdate="2014-01-01" gender="F" lastname="Wittlief" firstname="Isabelle" license="0">
              <RESULTS>
                <RESULT resultid="51" eventid="5" status="DSQ" swimtime="00:01:25.50" lane="3" heatid="5002" comment="Falscher Start." />
                <RESULT resultid="52" eventid="8" swimtime="00:00:46.72" lane="7" heatid="8002" />
                <RESULT resultid="53" eventid="10" swimtime="00:00:38.36" lane="8" heatid="10002" />
                <RESULT resultid="54" eventid="13" swimtime="00:03:17.04" lane="2" heatid="13002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:37.29" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="19" birthdate="2005-01-01" gender="M" lastname="Kwauka" firstname="Kevin" license="0">
              <RESULTS>
                <RESULT resultid="55" eventid="1" swimtime="00:00:18.76" lane="5" heatid="1006" />
                <RESULT resultid="56" eventid="5" swimtime="00:00:48.68" lane="8" heatid="5018" />
                <RESULT resultid="57" eventid="10" swimtime="00:00:20.19" lane="1" heatid="10018" />
                <RESULT resultid="58" eventid="12" swimtime="00:00:46.94" lane="8" heatid="12005" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="20" birthdate="2005-01-01" gender="F" lastname="Eweleit" firstname="Laura" license="0">
              <RESULTS>
                <RESULT resultid="59" eventid="1" swimtime="00:00:19.10" lane="4" heatid="1006" />
                <RESULT resultid="60" eventid="5" swimtime="00:00:45.09" lane="4" heatid="5017" />
                <RESULT resultid="61" eventid="10" swimtime="00:00:21.05" lane="8" heatid="10018" />
                <RESULT resultid="62" eventid="13" swimtime="00:01:40.80" lane="5" heatid="13012">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:48.54" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="21" birthdate="2010-01-01" gender="F" lastname="Haupt" firstname="Lena" license="0">
              <RESULTS>
                <RESULT resultid="63" eventid="5" swimtime="00:00:53.86" lane="5" heatid="5013" />
                <RESULT resultid="64" eventid="10" swimtime="00:00:25.13" lane="5" heatid="10013" />
                <RESULT resultid="65" eventid="13" swimtime="00:02:02.59" lane="5" heatid="13010">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:00.53" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="22" birthdate="2010-01-01" gender="F" lastname="Driescher" firstname="Leni" license="0">
              <RESULTS>
                <RESULT resultid="66" eventid="3" swimtime="00:05:26.64" lane="4" heatid="3004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:15.04" />
                    <SPLIT distance="200" swimtime="00:02:41.42" />
                    <SPLIT distance="300" swimtime="00:04:09.11" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="67" eventid="5" swimtime="00:01:13.40" lane="2" heatid="5009" />
                <RESULT resultid="68" eventid="10" swimtime="00:00:31.20" lane="6" heatid="10009" />
                <RESULT resultid="69" eventid="13" swimtime="00:02:43.33" lane="2" heatid="13007">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:17.66" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="23" birthdate="2011-01-01" gender="F" lastname="Eweleit" firstname="Lenja" license="0">
              <RESULTS>
                <RESULT resultid="70" eventid="3" swimtime="00:04:39.68" lane="1" heatid="3007">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:07.67" />
                    <SPLIT distance="200" swimtime="00:02:20.62" />
                    <SPLIT distance="300" swimtime="00:03:33.05" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="71" eventid="5" swimtime="00:00:58.82" lane="3" heatid="5012" />
                <RESULT resultid="72" eventid="10" swimtime="00:00:25.91" lane="7" heatid="10012" />
                <RESULT resultid="73" eventid="13" swimtime="00:02:10.21" lane="3" heatid="13009">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:03.28" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="24" birthdate="2009-01-01" gender="M" lastname="Vogler" firstname="Lennard" license="0">
              <RESULTS>
                <RESULT resultid="74" eventid="5" swimtime="00:01:15.13" lane="7" heatid="5005" />
                <RESULT resultid="75" eventid="10" swimtime="00:00:33.69" lane="5" heatid="10004" />
                <RESULT resultid="76" eventid="13" swimtime="00:02:52.12" lane="4" heatid="13003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:21.46" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="25" birthdate="2005-01-01" gender="F" lastname="Reinbach" firstname="Lilly" license="0">
              <RESULTS>
                <RESULT resultid="77" eventid="1" swimtime="00:00:23.25" lane="7" heatid="1004" />
                <RESULT resultid="78" eventid="5" swimtime="00:00:52.59" lane="5" heatid="5015" />
                <RESULT resultid="79" eventid="10" swimtime="00:00:25.39" lane="8" heatid="10015" />
                <RESULT resultid="80" eventid="13" swimtime="00:01:57.41" lane="3" heatid="13011">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:58.22" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="26" birthdate="2012-01-01" gender="F" lastname="Jeschke" firstname="Mira" license="0">
              <RESULTS>
                <RESULT resultid="81" eventid="3" swimtime="00:05:30.91" lane="5" heatid="3004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:16.62" />
                    <SPLIT distance="200" swimtime="00:02:41.59" />
                    <SPLIT distance="300" swimtime="00:04:11.42" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="82" eventid="5" swimtime="00:01:07.23" lane="5" heatid="5009" />
                <RESULT resultid="83" eventid="8" swimtime="00:00:32.29" lane="2" heatid="8004" />
                <RESULT resultid="84" eventid="10" swimtime="00:00:33.53" lane="8" heatid="10008" />
                <RESULT resultid="85" eventid="13" swimtime="00:02:37.26" lane="6" heatid="13007">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:17.53" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="27" birthdate="2007-01-01" gender="F" lastname="Götz" firstname="Zoe" license="0">
              <RESULTS>
                <RESULT resultid="86" eventid="1" swimtime="00:00:21.15" lane="8" heatid="1005" />
                <RESULT resultid="87" eventid="5" swimtime="00:00:51.89" lane="2" heatid="5016" />
                <RESULT resultid="88" eventid="6" swimtime="00:04:41.54" lane="7" heatid="6001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:06.83" />
                    <SPLIT distance="200" swimtime="00:02:19.32" />
                    <SPLIT distance="300" swimtime="00:03:32.24" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="89" eventid="10" swimtime="00:00:23.02" lane="1" heatid="10016" />
                <RESULT resultid="90" eventid="12" swimtime="00:00:50.76" lane="2" heatid="12004" />
                <RESULT resultid="91" eventid="13" swimtime="00:02:08.54" lane="2" heatid="13011">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:00.94" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY number="1" gender="X" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="18" eventid="14" swimtime="00:02:16.79" lane="5" heatid="14003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:43.17" />
                    <SPLIT distance="200" swimtime="00:01:31.02" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="15" number="1" />
                    <RELAYPOSITION athleteid="19" number="2" />
                    <RELAYPOSITION athleteid="20" number="3" />
                    <RELAYPOSITION athleteid="27" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="2" gender="X" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="19" eventid="14" swimtime="00:02:40.45" lane="4" heatid="14002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:50.62" />
                    <SPLIT distance="200" swimtime="00:01:44.90" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="14" number="1" />
                    <RELAYPOSITION athleteid="10" number="2" />
                    <RELAYPOSITION athleteid="21" number="3" />
                    <RELAYPOSITION athleteid="23" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="3" gender="X" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="20" eventid="14" swimtime="00:03:08.48" lane="1" heatid="14002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:54.18" />
                    <SPLIT distance="200" swimtime="00:02:00.84" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="17" number="1" />
                    <RELAYPOSITION athleteid="26" number="2" />
                    <RELAYPOSITION athleteid="16" number="3" />
                    <RELAYPOSITION athleteid="24" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="4" gender="X" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="21" eventid="14" swimtime="00:03:22.14" lane="5" heatid="14001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:57.76" />
                    <SPLIT distance="200" swimtime="00:02:08.20" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="25" number="1" />
                    <RELAYPOSITION athleteid="12" number="2" />
                    <RELAYPOSITION athleteid="22" number="3" />
                    <RELAYPOSITION athleteid="18" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB name="Tc submarin Pößneck" nation="GER" region="35" code="174116000">
          <ATHLETES>
            <ATHLETE athleteid="41" birthdate="2015-01-01" gender="F" lastname="Knoblich" firstname="Anna" license="0">
              <RESULTS>
                <RESULT resultid="123" eventid="2" swimtime="00:00:45.55" lane="7" heatid="2002" />
                <RESULT resultid="124" eventid="7" swimtime="00:00:49.79" lane="4" heatid="7001" />
                <RESULT resultid="125" eventid="11" swimtime="00:00:48.38" lane="2" heatid="11001" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="42" birthdate="2011-01-01" gender="M" lastname="Rattke" firstname="Carlos" license="0">
              <RESULTS>
                <RESULT resultid="126" eventid="3" swimtime="00:05:39.35" lane="7" heatid="3004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:18.37" />
                    <SPLIT distance="200" swimtime="00:02:48.18" />
                    <SPLIT distance="300" swimtime="00:04:19.41" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="127" eventid="5" swimtime="00:01:14.16" lane="6" heatid="5007" />
                <RESULT resultid="128" eventid="10" swimtime="00:00:33.92" lane="6" heatid="10007" />
                <RESULT resultid="129" eventid="12" swimtime="00:01:31.57" lane="1" heatid="12001" />
                <RESULT resultid="130" eventid="13" swimtime="00:02:37.72" lane="3" heatid="13006">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:18.66" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="44" birthdate="2007-01-01" gender="F" lastname="Näther" firstname="Emilia" license="0">
              <RESULTS>
                <RESULT resultid="136" eventid="1" swimtime="00:00:18.97" lane="6" heatid="1006" />
                <RESULT resultid="137" eventid="5" swimtime="00:00:46.63" lane="6" heatid="5017" />
                <RESULT resultid="138" eventid="10" swimtime="00:00:21.31" lane="2" heatid="10017" />
                <RESULT resultid="139" eventid="12" swimtime="00:00:48.58" lane="5" heatid="12004" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="45" birthdate="2013-01-01" gender="F" lastname="Dietzel" firstname="Hanna" license="0">
              <RESULTS>
                <RESULT resultid="140" eventid="5" swimtime="00:01:27.74" lane="1" heatid="5003" />
                <RESULT resultid="141" eventid="8" swimtime="00:00:42.23" lane="6" heatid="8001" />
                <RESULT resultid="142" eventid="10" swimtime="00:00:37.02" lane="8" heatid="10003" />
                <RESULT resultid="143" eventid="13" swimtime="00:03:14.60" lane="7" heatid="13002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:33.46" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="46" birthdate="2015-01-01" gender="F" lastname="Huber" firstname="Karla" license="0">
              <RESULTS>
                <RESULT resultid="144" eventid="2" swimtime="00:00:36.44" lane="6" heatid="2002" />
                <RESULT resultid="145" eventid="4" swimtime="00:00:18.34" lane="2" heatid="4001" />
                <RESULT resultid="146" eventid="7" swimtime="00:00:37.93" lane="2" heatid="7002" />
                <RESULT resultid="147" eventid="11" swimtime="00:00:44.45" lane="6" heatid="11001" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="47" birthdate="2014-01-01" gender="F" lastname="Cislak" firstname="Leni" license="0">
              <RESULTS>
                <RESULT resultid="148" eventid="5" swimtime="00:01:29.85" lane="4" heatid="5001" />
                <RESULT resultid="149" eventid="8" swimtime="00:00:44.94" lane="3" heatid="8001" />
                <RESULT resultid="150" eventid="10" swimtime="00:00:39.76" lane="4" heatid="10001" />
                <RESULT resultid="151" eventid="13" swimtime="00:03:27.21" lane="1" heatid="13003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:37.64" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="48" birthdate="2012-01-01" gender="F" lastname="Kraus" firstname="Letizia Marie" license="0">
              <RESULTS>
                <RESULT resultid="152" eventid="3" swimtime="00:04:31.68" lane="7" heatid="3007">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:01.95" />
                    <SPLIT distance="200" swimtime="00:02:12.09" />
                    <SPLIT distance="300" swimtime="00:03:23.94" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="153" eventid="5" swimtime="00:00:58.12" lane="8" heatid="5012" />
                <RESULT resultid="154" eventid="8" swimtime="00:00:29.34" lane="5" heatid="8004" />
                <RESULT resultid="155" eventid="10" swimtime="00:00:24.78" lane="8" heatid="10011" />
                <RESULT resultid="156" eventid="13" swimtime="00:02:06.62" lane="8" heatid="13009">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:00.65" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="49" birthdate="2016-01-01" gender="M" lastname="Kraus" firstname="Luan" license="0">
              <RESULTS>
                <RESULT resultid="157" eventid="2" swimtime="00:00:40.87" lane="5" heatid="2002" />
                <RESULT resultid="158" eventid="7" swimtime="00:00:40.59" lane="7" heatid="7002" />
                <RESULT resultid="159" eventid="11" swimtime="00:00:50.63" lane="7" heatid="11001" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="50" birthdate="2013-01-01" gender="F" lastname="Trunk" firstname="Mila" license="0">
              <RESULTS>
                <RESULT resultid="160" eventid="3" swimtime="00:05:47.10" lane="7" heatid="3003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:24.17" />
                    <SPLIT distance="200" swimtime="00:02:56.97" />
                    <SPLIT distance="300" swimtime="00:04:27.24" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="161" eventid="5" swimtime="00:01:12.77" lane="3" heatid="5005" />
                <RESULT resultid="162" eventid="8" swimtime="00:00:41.12" lane="3" heatid="8002" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="51" birthdate="2011-01-01" gender="M" lastname="Knoblich" firstname="Paul" license="0">
              <RESULTS>
                <RESULT resultid="163" eventid="3" swimtime="00:05:30.66" lane="6" heatid="3004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:17.32" />
                    <SPLIT distance="200" swimtime="00:02:46.38" />
                    <SPLIT distance="300" swimtime="00:04:15.59" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="164" eventid="5" swimtime="00:01:07.19" lane="4" heatid="5008" />
                <RESULT resultid="165" eventid="10" swimtime="00:00:32.48" lane="7" heatid="10007" />
                <RESULT resultid="166" eventid="12" swimtime="00:01:25.54" lane="7" heatid="12001" />
                <RESULT resultid="167" eventid="13" swimtime="00:02:37.36" lane="4" heatid="13006">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:18.98" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="52" birthdate="2013-01-01" gender="F" lastname="Huber" firstname="Sina" license="0">
              <RESULTS>
                <RESULT resultid="168" eventid="3" swimtime="00:05:49.49" lane="4" heatid="3003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:25.06" />
                    <SPLIT distance="200" swimtime="00:02:56.16" />
                    <SPLIT distance="300" swimtime="00:04:26.24" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="169" eventid="5" swimtime="00:01:14.67" lane="8" heatid="5006" />
                <RESULT resultid="170" eventid="8" swimtime="00:00:35.38" lane="8" heatid="8003" />
                <RESULT resultid="171" eventid="10" swimtime="00:00:32.55" lane="2" heatid="10006" />
                <RESULT resultid="172" eventid="13" swimtime="00:02:49.88" lane="1" heatid="13006">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:23.64" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="53" birthdate="2010-01-01" gender="F" lastname="Matthes" firstname="Sophie" license="0">
              <RESULTS>
                <RESULT resultid="173" eventid="3" swimtime="00:05:10.51" lane="8" heatid="3005">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:13.49" />
                    <SPLIT distance="200" swimtime="00:02:37.25" />
                    <SPLIT distance="300" swimtime="00:04:00.26" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="174" eventid="5" swimtime="00:01:03.36" lane="5" heatid="5012" />
                <RESULT resultid="175" eventid="10" swimtime="00:00:27.40" lane="6" heatid="10012" />
                <RESULT resultid="176" eventid="12" swimtime="00:01:02.56" lane="2" heatid="12003" />
                <RESULT resultid="177" eventid="13" status="DSQ" swimtime="00:02:33.06" lane="7" heatid="13008" comment="Tauchzüge außerhalb der 15m-Zone bei ca. 125 Meter.">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:16.91" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="55" birthdate="2013-01-01" gender="F" lastname="Schmidt" firstname="Ylva" license="0">
              <RESULTS>
                <RESULT resultid="179" eventid="3" swimtime="00:06:03.87" lane="6" heatid="3002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:24.04" />
                    <SPLIT distance="200" swimtime="00:02:59.04" />
                    <SPLIT distance="300" swimtime="00:04:34.21" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="180" eventid="5" swimtime="00:01:13.95" lane="1" heatid="5005" />
                <RESULT resultid="181" eventid="8" swimtime="00:00:34.71" lane="4" heatid="8003" />
                <RESULT resultid="182" eventid="10" swimtime="00:00:33.18" lane="1" heatid="10006" />
                <RESULT resultid="183" eventid="13" swimtime="00:02:56.77" lane="4" heatid="13004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:28.10" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="56" birthdate="2013-01-01" gender="F" lastname="Werner" firstname="Zoe" license="0">
              <RESULTS>
                <RESULT resultid="184" eventid="3" swimtime="00:05:48.05" lane="5" heatid="3003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:23.75" />
                    <SPLIT distance="200" swimtime="00:02:56.31" />
                    <SPLIT distance="300" swimtime="00:04:26.63" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="185" eventid="5" swimtime="00:01:17.25" lane="8" heatid="5005" />
                <RESULT resultid="186" eventid="8" swimtime="00:00:37.11" lane="6" heatid="8002" />
                <RESULT resultid="187" eventid="10" swimtime="00:00:35.74" lane="2" heatid="10004" />
                <RESULT resultid="188" eventid="13" swimtime="00:02:52.36" lane="1" heatid="13005">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:26.24" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="TSC Rostock 1957 e.V." nation="GER" region="22" code="0">
          <ATHLETES>
            <ATHLETE athleteid="104" birthdate="2010-01-01" gender="F" lastname="Timmer" firstname="Anna Fee" license="0">
              <RESULTS>
                <RESULT resultid="331" eventid="5" swimtime="00:01:06.53" lane="4" heatid="5009" />
                <RESULT resultid="332" eventid="10" swimtime="00:00:29.61" lane="3" heatid="10008" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="105" birthdate="2009-01-01" gender="F" lastname="Mende" firstname="Carla" license="0">
              <RESULTS>
                <RESULT resultid="333" eventid="1" swimtime="00:00:25.95" lane="1" heatid="1002" />
                <RESULT resultid="334" eventid="5" swimtime="00:01:05.66" lane="5" heatid="5010" />
                <RESULT resultid="335" eventid="12" swimtime="00:01:03.36" lane="3" heatid="12002" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="106" birthdate="2011-01-01" gender="F" lastname="Drews" firstname="Elsa" license="0">
              <RESULTS>
                <RESULT resultid="336" eventid="5" swimtime="00:01:11.84" lane="2" heatid="5007" />
                <RESULT resultid="337" eventid="10" swimtime="00:00:31.40" lane="6" heatid="10008" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="107" birthdate="2010-01-01" gender="F" lastname="Buch" firstname="Freya" license="0">
              <RESULTS>
                <RESULT resultid="338" eventid="3" swimtime="00:04:44.28" lane="6" heatid="3007">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:05.96" />
                    <SPLIT distance="200" swimtime="00:02:20.16" />
                    <SPLIT distance="300" swimtime="00:03:35.02" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="339" eventid="5" swimtime="00:01:00.12" lane="6" heatid="5011" />
                <RESULT resultid="340" eventid="6" status="DNS" swimtime="00:00:00.00" lane="1" heatid="6001" />
                <RESULT resultid="341" eventid="12" swimtime="00:01:04.69" lane="4" heatid="12002" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="108" birthdate="2011-01-01" gender="M" lastname="Behrend" firstname="Gustav" license="0">
              <RESULTS>
                <RESULT resultid="342" eventid="10" swimtime="00:00:31.85" lane="7" heatid="10009" />
                <RESULT resultid="343" eventid="12" swimtime="00:01:22.75" lane="5" heatid="12001" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="109" birthdate="2011-01-01" gender="F" lastname="Beerbaum" firstname="Isabella" license="0">
              <RESULTS>
                <RESULT resultid="344" eventid="5" swimtime="00:01:08.74" lane="1" heatid="5009" />
                <RESULT resultid="345" eventid="10" swimtime="00:00:30.29" lane="5" heatid="10008" />
                <RESULT resultid="346" eventid="12" swimtime="00:01:18.29" lane="3" heatid="12001" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="110" birthdate="2009-01-01" gender="M" lastname="Wippler" firstname="Jannik" license="0">
              <RESULTS>
                <RESULT resultid="347" eventid="1" swimtime="00:00:29.29" lane="5" heatid="1001" />
                <RESULT resultid="348" eventid="3" swimtime="00:05:00.56" lane="3" heatid="3005">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:09.70" />
                    <SPLIT distance="200" swimtime="00:02:28.97" />
                    <SPLIT distance="300" swimtime="00:03:48.32" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="349" eventid="5" swimtime="00:01:02.57" lane="6" heatid="5010" />
                <RESULT resultid="350" eventid="12" swimtime="00:01:14.99" lane="7" heatid="12002" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="111" birthdate="2010-01-01" gender="F" lastname="Reichardt" firstname="Jula" license="0">
              <RESULTS>
                <RESULT resultid="351" eventid="3" swimtime="00:04:47.49" lane="6" heatid="3006">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:05.07" />
                    <SPLIT distance="200" swimtime="00:02:22.02" />
                    <SPLIT distance="300" swimtime="00:03:38.40" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="352" eventid="5" swimtime="00:01:00.24" lane="3" heatid="5011" />
                <RESULT resultid="353" eventid="10" swimtime="00:00:27.37" lane="4" heatid="10010" />
                <RESULT resultid="354" eventid="12" swimtime="00:01:04.47" lane="6" heatid="12002" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="112" birthdate="2010-01-01" gender="M" lastname="Koslov" firstname="Luis" license="0">
              <RESULTS>
                <RESULT resultid="355" eventid="3" swimtime="00:04:40.98" lane="4" heatid="3006">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:04.54" />
                    <SPLIT distance="200" swimtime="00:02:18.50" />
                    <SPLIT distance="300" swimtime="00:03:32.26" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="356" eventid="5" swimtime="00:00:57.77" lane="7" heatid="5003" />
                <RESULT resultid="357" eventid="6" status="DNS" swimtime="00:00:00.00" lane="8" heatid="6001" />
                <RESULT resultid="358" eventid="10" swimtime="00:00:26.34" lane="3" heatid="10012" />
                <RESULT resultid="359" eventid="12" swimtime="00:00:58.33" lane="1" heatid="12003" />
                <RESULT resultid="360" eventid="13" swimtime="00:02:13.44" lane="7" heatid="13009">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:04.85" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="113" birthdate="2010-01-01" gender="F" lastname="Peetz" firstname="Marthe" license="0">
              <RESULTS>
                <RESULT resultid="361" eventid="5" status="DSQ" swimtime="00:01:10.85" lane="6" heatid="5009" comment="flascher Start" />
                <RESULT resultid="362" eventid="10" swimtime="00:00:30.54" lane="1" heatid="10009" />
                <RESULT resultid="363" eventid="12" swimtime="00:01:13.62" lane="6" heatid="12001" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY number="1" gender="X" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="364" eventid="14" swimtime="00:03:08.69" lane="6" heatid="14002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:59.06" />
                    <SPLIT distance="200" swimtime="00:02:04.58" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="110" number="1" />
                    <RELAYPOSITION athleteid="107" number="2" />
                    <RELAYPOSITION athleteid="113" number="3" />
                    <RELAYPOSITION athleteid="111" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" gender="X" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="365" eventid="14" swimtime="00:03:09.57" lane="2" heatid="14002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:59.65" />
                    <SPLIT distance="200" swimtime="00:02:06.99" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="105" number="1" />
                    <RELAYPOSITION athleteid="112" number="2" />
                    <RELAYPOSITION athleteid="104" number="3" />
                    <RELAYPOSITION athleteid="106" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB name="TSC Schwandorf e.V." nation="GER" region="34" code="0">
          <ATHLETES>
            <ATHLETE athleteid="57" birthdate="2004-01-01" gender="F" lastname="Kohler" firstname="Nina" license="0">
              <RESULTS>
                <RESULT resultid="189" eventid="1" swimtime="00:00:18.28" lane="1" heatid="1007" />
                <RESULT resultid="190" eventid="5" swimtime="00:00:44.41" lane="1" heatid="5018" />
                <RESULT resultid="191" eventid="10" swimtime="00:00:19.99" lane="4" heatid="10017" />
                <RESULT resultid="192" eventid="12" swimtime="00:00:42.47" lane="3" heatid="12005" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="TSG TU Ilmenau 56 e.V." nation="GER" region="35" code="0">
          <ATHLETES>
            <ATHLETE athleteid="163" birthdate="2001-01-01" gender="M" lastname="Pohl" firstname="Enrico" license="0">
              <RESULTS>
                <RESULT resultid="537" eventid="1" swimtime="00:00:15.95" lane="4" heatid="1007" />
                <RESULT resultid="538" eventid="5" swimtime="00:00:38.79" lane="4" heatid="5018" />
                <RESULT resultid="539" eventid="10" swimtime="00:00:17.42" lane="4" heatid="10018" />
                <RESULT resultid="540" eventid="12" swimtime="00:00:39.38" lane="4" heatid="12005" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="164" birthdate="2013-01-01" gender="M" lastname="Albrecht" firstname="Leopold" license="0">
              <RESULTS>
                <RESULT resultid="541" eventid="5" swimtime="00:01:18.99" lane="5" heatid="5001" />
                <RESULT resultid="542" eventid="8" swimtime="00:00:47.47" lane="7" heatid="8001" />
                <RESULT resultid="543" eventid="10" swimtime="00:00:36.43" lane="2" heatid="10001" />
                <RESULT resultid="544" eventid="13" swimtime="00:02:57.85" lane="5" heatid="13001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:30.22" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="165" birthdate="2008-01-01" gender="F" lastname="Liebhold" firstname="Lotta" license="0">
              <RESULTS>
                <RESULT resultid="545" eventid="1" swimtime="00:00:24.68" lane="6" heatid="1002" />
                <RESULT resultid="546" eventid="3" swimtime="00:04:45.04" lane="4" heatid="3007">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:05.71" />
                    <SPLIT distance="200" swimtime="00:02:19.80" />
                    <SPLIT distance="300" swimtime="00:03:35.00" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="547" eventid="5" swimtime="00:00:56.45" lane="8" heatid="5013" />
                <RESULT resultid="548" eventid="10" swimtime="00:00:25.13" lane="5" heatid="10012" />
                <RESULT resultid="549" eventid="12" swimtime="00:00:59.88" lane="5" heatid="12002" />
                <RESULT resultid="550" eventid="13" swimtime="00:02:11.75" lane="4" heatid="13009">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:04.04" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="166" birthdate="2007-01-01" gender="M" lastname="Stuwe" firstname="Paul" license="0">
              <RESULTS>
                <RESULT resultid="551" eventid="1" swimtime="00:00:20.97" lane="5" heatid="1004" />
                <RESULT resultid="552" eventid="3" swimtime="00:04:20.99" lane="8" heatid="3009">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:59.93" />
                    <SPLIT distance="200" swimtime="00:02:05.86" />
                    <SPLIT distance="300" swimtime="00:03:13.19" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="553" eventid="6" swimtime="00:04:19.19" lane="3" heatid="6001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:55.99" />
                    <SPLIT distance="200" swimtime="00:02:02.29" />
                    <SPLIT distance="300" swimtime="00:03:10.35" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="554" eventid="10" swimtime="00:00:23.19" lane="4" heatid="10014" />
                <RESULT resultid="555" eventid="13" swimtime="00:01:57.16" lane="6" heatid="13009">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:55.67" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="167" birthdate="2016-01-01" gender="M" lastname="Stuwe" firstname="Piet" license="0">
              <RESULTS>
                <RESULT resultid="556" eventid="2" swimtime="00:00:50.22" lane="8" heatid="2002" />
                <RESULT resultid="557" eventid="7" swimtime="00:00:56.80" lane="5" heatid="7001" />
                <RESULT resultid="558" eventid="11" swimtime="00:00:48.07" lane="1" heatid="11001" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
      </CLUBS>
    </MEET>
  </MEETS>
</LENEX>
