<?xml version="1.0" encoding="UTF-8"?>
<LENEX version="3.0">
  <CONSTRUCTOR name="EasyWk" version="5.23 BETA" registration="">
    <CONTACT name="Bjoern Stickan" internet="http://www.easywk.de" email="info@easywk.de" />
  </CONSTRUCTOR>
  <MEETS>
    <MEET city="Erfurt" course="LCM" name="Fühlingspokal und 42. Offene Süddeutsche Meisterschaften im Finswimming" nation="GER" organizer="Tauchsportclub Erfurt e.V." hostclub="LTV Baden, Bayern, Hessen Rheinland-Pfalz, Saarland, Thüringen, Würtemberg" deadline="2023-03-15" timing="AUTOMATIC">
      <CONTACT city="Erfurt" email="sdm@fs-ergebnisse.de" internet="www.fs-ergebnisse.de/2023/sdm" name="Sabine Delcuvé, Meldeservice SDM 2023" phone="0160 99161353" />
      <AGEDATE type="YEAR" value="2023-01-01" />
      <SESSIONS>
        <SESSION number="1" date="2023-03-25" daytime="10:20" officialmeeting="09:30" warmupfrom="09:00">
          <EVENTS>
            <EVENT eventid="1" number="1" gender="F" round="TIM">
              <SWIMSTYLE stroke="SURFACE" relaycount="1" distance="100" />
              <FEE value="500" currency="EUR" />
              <HEATS>
                <HEAT heatid="1001" number="1" />
                <HEAT heatid="1002" number="2" />
                <HEAT heatid="1003" number="3" />
                <HEAT heatid="1004" number="4" />
                <HEAT heatid="1005" number="5" />
                <HEAT heatid="1006" number="6" />
                <HEAT heatid="1007" number="7" />
                <HEAT heatid="1008" number="8" />
                <HEAT heatid="1009" number="9" />
                <HEAT heatid="1010" number="10" />
                <HEAT heatid="1011" number="11" />
                <HEAT heatid="1012" number="12" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="4" agemax="9" agemin="3" name="Jahrgang 2014 und jünger - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="3" resultid="184" />
                    <RANKING place="1" resultid="294" />
                    <RANKING place="4" resultid="423" />
                    <RANKING place="2" resultid="705" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="10" agemin="10" name="Jahrgang 2013 - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="5" resultid="293" />
                    <RANKING place="6" resultid="431" />
                    <RANKING place="1" resultid="1004" />
                    <RANKING place="4" resultid="1005" />
                    <RANKING place="2" resultid="1006" />
                    <RANKING place="3" resultid="1008" />
                    <RANKING place="7" resultid="1009" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6" agemax="11" agemin="11" name="Jahrgang 2012 - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="3" resultid="181" />
                    <RANKING place="1" resultid="182" />
                    <RANKING place="10" resultid="430" />
                    <RANKING place="7" resultid="432" />
                    <RANKING place="5" resultid="702" />
                    <RANKING place="9" resultid="793" />
                    <RANKING place="4" resultid="794" />
                    <RANKING place="8" resultid="795" />
                    <RANKING place="6" resultid="798" />
                    <RANKING place="2" resultid="1002" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7" agemax="12" agemin="12" name="Jahrgang 2011 - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="2" resultid="125" />
                    <RANKING place="3" resultid="183" />
                    <RANKING place="6" resultid="290" />
                    <RANKING place="9" resultid="291" />
                    <RANKING place="7" resultid="292" />
                    <RANKING place="5" resultid="429" />
                    <RANKING place="8" resultid="704" />
                    <RANKING place="1" resultid="791" />
                    <RANKING place="4" resultid="1003" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8" agemax="13" agemin="13" name="Jahrgang 2010 - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="2" resultid="124" />
                    <RANKING place="5" resultid="427" />
                    <RANKING place="6" resultid="428" />
                    <RANKING place="4" resultid="701" />
                    <RANKING place="7" resultid="703" />
                    <RANKING place="1" resultid="786" />
                    <RANKING place="8" resultid="797" />
                    <RANKING place="3" resultid="1001" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9" agemax="14" agemin="14" name="Jahrgang 2009 - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="7" resultid="63" />
                    <RANKING place="2" resultid="176" />
                    <RANKING place="5" resultid="180" />
                    <RANKING place="3" resultid="289" />
                    <RANKING place="4" resultid="668" />
                    <RANKING place="8" resultid="669" />
                    <RANKING place="1" resultid="783" />
                    <RANKING place="6" resultid="792" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10" agemax="15" agemin="15" name="Jahrgang 2008 - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="1" resultid="178" />
                    <RANKING place="2" resultid="698" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11" agemax="16" agemin="16" name="Jahrgang 2007 - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="5" resultid="5" />
                    <RANKING place="3" resultid="62" />
                    <RANKING place="4" resultid="126" />
                    <RANKING place="1" resultid="146" />
                    <RANKING place="2" resultid="999" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="12" agemax="17" agemin="17" name="Jahrgang 2006 - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="1" resultid="287" />
                    <RANKING place="2" resultid="288" />
                    <RANKING place="4" resultid="667" />
                    <RANKING place="5" resultid="699" />
                    <RANKING place="3" resultid="785" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="13" agemax="21" agemin="18" name="Juniorinnen - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="1" resultid="122" />
                    <RANKING place="4" resultid="175" />
                    <RANKING place="2" resultid="286" />
                    <RANKING place="7" resultid="424" />
                    <RANKING place="5" resultid="425" />
                    <RANKING place="8" resultid="787" />
                    <RANKING place="3" resultid="998" />
                    <RANKING place="6" resultid="1000" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="14" agemax="28" agemin="3" name="Offene Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="22" resultid="4" />
                    <RANKING place="52" resultid="5" />
                    <RANKING place="20" resultid="62" />
                    <RANKING place="44" resultid="63" />
                    <RANKING place="1" resultid="122" />
                    <RANKING place="30" resultid="124" />
                    <RANKING place="39" resultid="125" />
                    <RANKING place="48" resultid="126" />
                    <RANKING place="7" resultid="146" />
                    <RANKING place="4" resultid="148" />
                    <RANKING place="3" resultid="149" />
                    <RANKING place="6" resultid="175" />
                    <RANKING place="16" resultid="176" />
                    <RANKING place="21" resultid="177" />
                    <RANKING place="15" resultid="178" />
                    <RANKING place="29" resultid="180" />
                    <RANKING place="35" resultid="181" />
                    <RANKING place="31" resultid="182" />
                    <RANKING place="41" resultid="183" />
                    <RANKING place="70" resultid="184" />
                    <RANKING place="2" resultid="286" />
                    <RANKING place="10" resultid="287" />
                    <RANKING place="17" resultid="288" />
                    <RANKING place="23" resultid="289" />
                    <RANKING place="49" resultid="290" />
                    <RANKING place="62" resultid="291" />
                    <RANKING place="53" resultid="292" />
                    <RANKING place="64" resultid="293" />
                    <RANKING place="68" resultid="294" />
                    <RANKING place="71" resultid="423" />
                    <RANKING place="12" resultid="424" />
                    <RANKING place="8" resultid="425" />
                    <RANKING place="37" resultid="427" />
                    <RANKING place="42" resultid="428" />
                    <RANKING place="46" resultid="429" />
                    <RANKING place="67" resultid="430" />
                    <RANKING place="65" resultid="431" />
                    <RANKING place="54" resultid="432" />
                    <RANKING place="24" resultid="667" />
                    <RANKING place="25" resultid="668" />
                    <RANKING place="50" resultid="669" />
                    <RANKING place="18" resultid="697" />
                    <RANKING place="28" resultid="698" />
                    <RANKING place="27" resultid="699" />
                    <RANKING place="36" resultid="701" />
                    <RANKING place="47" resultid="702" />
                    <RANKING place="45" resultid="703" />
                    <RANKING place="58" resultid="704" />
                    <RANKING place="69" resultid="705" />
                    <RANKING place="9" resultid="783" />
                    <RANKING place="19" resultid="785" />
                    <RANKING place="14" resultid="786" />
                    <RANKING place="26" resultid="787" />
                    <RANKING place="38" resultid="791" />
                    <RANKING place="33" resultid="792" />
                    <RANKING place="56" resultid="793" />
                    <RANKING place="40" resultid="794" />
                    <RANKING place="55" resultid="795" />
                    <RANKING place="63" resultid="797" />
                    <RANKING place="51" resultid="798" />
                    <RANKING place="5" resultid="998" />
                    <RANKING place="13" resultid="999" />
                    <RANKING place="11" resultid="1000" />
                    <RANKING place="34" resultid="1001" />
                    <RANKING place="32" resultid="1002" />
                    <RANKING place="43" resultid="1003" />
                    <RANKING place="57" resultid="1004" />
                    <RANKING place="61" resultid="1005" />
                    <RANKING place="59" resultid="1006" />
                    <RANKING place="60" resultid="1008" />
                    <RANKING place="66" resultid="1009" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="19" agemax="28" agemin="3" name="Offene internationale Wertung">
                  <RANKINGS>
                    <RANKING place="25" resultid="4" />
                    <RANKING place="60" resultid="5" />
                    <RANKING place="23" resultid="62" />
                    <RANKING place="52" resultid="63" />
                    <RANKING place="12" resultid="73" />
                    <RANKING place="18" resultid="75" />
                    <RANKING place="36" resultid="76" />
                    <RANKING place="1" resultid="122" />
                    <RANKING place="35" resultid="124" />
                    <RANKING place="47" resultid="125" />
                    <RANKING place="56" resultid="126" />
                    <RANKING place="7" resultid="146" />
                    <RANKING place="4" resultid="148" />
                    <RANKING place="3" resultid="149" />
                    <RANKING place="6" resultid="175" />
                    <RANKING place="19" resultid="176" />
                    <RANKING place="24" resultid="177" />
                    <RANKING place="17" resultid="178" />
                    <RANKING place="34" resultid="180" />
                    <RANKING place="42" resultid="181" />
                    <RANKING place="37" resultid="182" />
                    <RANKING place="49" resultid="183" />
                    <RANKING place="78" resultid="184" />
                    <RANKING place="2" resultid="286" />
                    <RANKING place="10" resultid="287" />
                    <RANKING place="20" resultid="288" />
                    <RANKING place="26" resultid="289" />
                    <RANKING place="57" resultid="290" />
                    <RANKING place="70" resultid="291" />
                    <RANKING place="61" resultid="292" />
                    <RANKING place="72" resultid="293" />
                    <RANKING place="76" resultid="294" />
                    <RANKING place="15" resultid="381" />
                    <RANKING place="27" resultid="382" />
                    <RANKING place="33" resultid="383" />
                    <RANKING place="40" resultid="384" />
                    <RANKING place="79" resultid="423" />
                    <RANKING place="13" resultid="424" />
                    <RANKING place="8" resultid="425" />
                    <RANKING place="44" resultid="427" />
                    <RANKING place="50" resultid="428" />
                    <RANKING place="54" resultid="429" />
                    <RANKING place="75" resultid="430" />
                    <RANKING place="73" resultid="431" />
                    <RANKING place="62" resultid="432" />
                    <RANKING place="45" resultid="658" />
                    <RANKING place="28" resultid="667" />
                    <RANKING place="29" resultid="668" />
                    <RANKING place="58" resultid="669" />
                    <RANKING place="21" resultid="697" />
                    <RANKING place="32" resultid="698" />
                    <RANKING place="31" resultid="699" />
                    <RANKING place="43" resultid="701" />
                    <RANKING place="55" resultid="702" />
                    <RANKING place="53" resultid="703" />
                    <RANKING place="66" resultid="704" />
                    <RANKING place="77" resultid="705" />
                    <RANKING place="9" resultid="783" />
                    <RANKING place="22" resultid="785" />
                    <RANKING place="16" resultid="786" />
                    <RANKING place="30" resultid="787" />
                    <RANKING place="46" resultid="791" />
                    <RANKING place="39" resultid="792" />
                    <RANKING place="64" resultid="793" />
                    <RANKING place="48" resultid="794" />
                    <RANKING place="63" resultid="795" />
                    <RANKING place="71" resultid="797" />
                    <RANKING place="59" resultid="798" />
                    <RANKING place="5" resultid="998" />
                    <RANKING place="14" resultid="999" />
                    <RANKING place="11" resultid="1000" />
                    <RANKING place="41" resultid="1001" />
                    <RANKING place="38" resultid="1002" />
                    <RANKING place="51" resultid="1003" />
                    <RANKING place="65" resultid="1004" />
                    <RANKING place="69" resultid="1005" />
                    <RANKING place="67" resultid="1006" />
                    <RANKING place="68" resultid="1008" />
                    <RANKING place="74" resultid="1009" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15" agemax="44" agemin="29" name="Master A - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="1" resultid="788" />
                    <RANKING place="3" resultid="789" />
                    <RANKING place="2" resultid="958" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="16" agemax="54" agemin="45" name="Master B - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="1" resultid="426" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="17" agemax="-1" agemin="55" name="Master C - Süddeutsche Wertung" />
                <AGEGROUP agegroupid="18" agemax="-1" agemin="29" name="Offene internationale Wertung Master">
                  <RANKINGS>
                    <RANKING place="1" resultid="426" />
                    <RANKING place="2" resultid="788" />
                    <RANKING place="4" resultid="789" />
                    <RANKING place="3" resultid="958" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="2" number="2" gender="M" round="TIM">
              <SWIMSTYLE stroke="SURFACE" relaycount="1" distance="100" />
              <FEE value="500" currency="EUR" />
              <HEATS>
                <HEAT heatid="2001" number="1" />
                <HEAT heatid="2002" number="2" />
                <HEAT heatid="2003" number="3" />
                <HEAT heatid="2004" number="4" />
                <HEAT heatid="2005" number="5" />
                <HEAT heatid="2006" number="6" />
                <HEAT heatid="2007" number="7" />
                <HEAT heatid="2008" number="8" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="4" agemax="9" agemin="3" name="Jahrgang 2014 und jünger - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="2" resultid="12" />
                    <RANKING place="1" resultid="300" />
                    <RANKING place="3" resultid="443" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="10" agemin="10" name="Jahrgang 2013 - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="2" resultid="11" />
                    <RANKING place="1" resultid="191" />
                    <RANKING place="3" resultid="192" />
                    <RANKING place="4" resultid="1012" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6" agemax="11" agemin="11" name="Jahrgang 2012 - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="1" resultid="190" />
                    <RANKING place="2" resultid="299" />
                    <RANKING place="3" resultid="671" />
                    <RANKING place="4" resultid="807" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7" agemax="12" agemin="12" name="Jahrgang 2011 - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="2" resultid="189" />
                    <RANKING place="3" resultid="298" />
                    <RANKING place="1" resultid="438" />
                    <RANKING place="6" resultid="708" />
                    <RANKING place="7" resultid="709" />
                    <RANKING place="5" resultid="1010" />
                    <RANKING place="4" resultid="1011" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8" agemax="13" agemin="13" name="Jahrgang 2010 - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="2" resultid="439" />
                    <RANKING place="1" resultid="802" />
                    <RANKING place="3" resultid="804" />
                    <RANKING place="4" resultid="806" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9" agemax="14" agemin="14" name="Jahrgang 2009 - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="2" resultid="8" />
                    <RANKING place="3" resultid="9" />
                    <RANKING place="1" resultid="297" />
                    <RANKING place="4" resultid="441" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10" agemax="15" agemin="15" name="Jahrgang 2008 - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="3" resultid="7" />
                    <RANKING place="1" resultid="295" />
                    <RANKING place="2" resultid="801" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11" agemax="16" agemin="16" name="Jahrgang 2007 - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="1" resultid="707" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="12" agemax="17" agemin="17" name="Jahrgang 2006 - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="3" resultid="6" />
                    <RANKING place="2" resultid="435" />
                    <RANKING place="1" resultid="799" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="13" agemax="21" agemin="18" name="Junioren - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="1" resultid="185" />
                    <RANKING place="5" resultid="188" />
                    <RANKING place="2" resultid="433" />
                    <RANKING place="3" resultid="434" />
                    <RANKING place="4" resultid="436" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="14" agemax="28" agemin="3" name="Offene Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="9" resultid="6" />
                    <RANKING place="11" resultid="7" />
                    <RANKING place="15" resultid="8" />
                    <RANKING place="20" resultid="9" />
                    <RANKING place="30" resultid="11" />
                    <RANKING place="38" resultid="12" />
                    <RANKING place="3" resultid="185" />
                    <RANKING place="13" resultid="188" />
                    <RANKING place="18" resultid="189" />
                    <RANKING place="24" resultid="190" />
                    <RANKING place="27" resultid="191" />
                    <RANKING place="34" resultid="192" />
                    <RANKING place="5" resultid="295" />
                    <RANKING place="14" resultid="297" />
                    <RANKING place="25" resultid="298" />
                    <RANKING place="31" resultid="299" />
                    <RANKING place="33" resultid="300" />
                    <RANKING place="4" resultid="433" />
                    <RANKING place="6" resultid="434" />
                    <RANKING place="7" resultid="435" />
                    <RANKING place="8" resultid="436" />
                    <RANKING place="17" resultid="438" />
                    <RANKING place="19" resultid="439" />
                    <RANKING place="23" resultid="441" />
                    <RANKING place="39" resultid="443" />
                    <RANKING place="32" resultid="671" />
                    <RANKING place="2" resultid="706" />
                    <RANKING place="12" resultid="707" />
                    <RANKING place="29" resultid="708" />
                    <RANKING place="37" resultid="709" />
                    <RANKING place="1" resultid="799" />
                    <RANKING place="9" resultid="801" />
                    <RANKING place="16" resultid="802" />
                    <RANKING place="21" resultid="804" />
                    <RANKING place="22" resultid="806" />
                    <RANKING place="35" resultid="807" />
                    <RANKING place="28" resultid="1010" />
                    <RANKING place="26" resultid="1011" />
                    <RANKING place="36" resultid="1012" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="19" agemax="28" agemin="3" name="Offene internationale Wertung">
                  <RANKINGS>
                    <RANKING place="14" resultid="6" />
                    <RANKING place="16" resultid="7" />
                    <RANKING place="20" resultid="8" />
                    <RANKING place="26" resultid="9" />
                    <RANKING place="36" resultid="11" />
                    <RANKING place="44" resultid="12" />
                    <RANKING place="1" resultid="77" />
                    <RANKING place="6" resultid="78" />
                    <RANKING place="13" resultid="79" />
                    <RANKING place="11" resultid="80" />
                    <RANKING place="5" resultid="185" />
                    <RANKING place="18" resultid="188" />
                    <RANKING place="24" resultid="189" />
                    <RANKING place="30" resultid="190" />
                    <RANKING place="33" resultid="191" />
                    <RANKING place="40" resultid="192" />
                    <RANKING place="8" resultid="295" />
                    <RANKING place="19" resultid="297" />
                    <RANKING place="31" resultid="298" />
                    <RANKING place="37" resultid="299" />
                    <RANKING place="39" resultid="300" />
                    <RANKING place="4" resultid="385" />
                    <RANKING place="21" resultid="386" />
                    <RANKING place="7" resultid="433" />
                    <RANKING place="9" resultid="434" />
                    <RANKING place="10" resultid="435" />
                    <RANKING place="12" resultid="436" />
                    <RANKING place="23" resultid="438" />
                    <RANKING place="25" resultid="439" />
                    <RANKING place="29" resultid="441" />
                    <RANKING place="45" resultid="443" />
                    <RANKING place="38" resultid="671" />
                    <RANKING place="3" resultid="706" />
                    <RANKING place="17" resultid="707" />
                    <RANKING place="35" resultid="708" />
                    <RANKING place="43" resultid="709" />
                    <RANKING place="2" resultid="799" />
                    <RANKING place="14" resultid="801" />
                    <RANKING place="22" resultid="802" />
                    <RANKING place="27" resultid="804" />
                    <RANKING place="28" resultid="806" />
                    <RANKING place="41" resultid="807" />
                    <RANKING place="34" resultid="1010" />
                    <RANKING place="32" resultid="1011" />
                    <RANKING place="42" resultid="1012" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15" agemax="44" agemin="29" name="Master A - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="1" resultid="150" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="16" agemax="54" agemin="45" name="Master B - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="2" resultid="296" />
                    <RANKING place="1" resultid="800" />
                    <RANKING place="3" resultid="803" />
                    <RANKING place="4" resultid="964" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="17" agemax="-1" agemin="55" name="Master C - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="1" resultid="118" />
                    <RANKING place="2" resultid="440" />
                    <RANKING place="3" resultid="442" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="18" agemax="-1" agemin="29" name="Offene internationale Wertung Master">
                  <RANKINGS>
                    <RANKING place="5" resultid="118" />
                    <RANKING place="2" resultid="150" />
                    <RANKING place="4" resultid="296" />
                    <RANKING place="8" resultid="440" />
                    <RANKING place="9" resultid="442" />
                    <RANKING place="3" resultid="800" />
                    <RANKING place="6" resultid="803" />
                    <RANKING place="1" resultid="953" />
                    <RANKING place="7" resultid="964" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="3" number="3" gender="F" round="TIM">
              <SWIMSTYLE stroke="BIFIN" relaycount="1" distance="100" />
              <FEE value="500" currency="EUR" />
              <HEATS>
                <HEAT heatid="3001" number="1" />
                <HEAT heatid="3002" number="2" />
                <HEAT heatid="3003" number="3" />
                <HEAT heatid="3004" number="4" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="4" agemax="9" agemin="3" name="Jahrgang 2014 und jünger - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="3" resultid="416" />
                    <RANKING place="5" resultid="990" />
                    <RANKING place="2" resultid="991" />
                    <RANKING place="1" resultid="992" />
                    <RANKING place="4" resultid="993" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="10" agemin="10" name="Jahrgang 2013 - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="3" resultid="281" />
                    <RANKING place="8" resultid="775" />
                    <RANKING place="5" resultid="776" />
                    <RANKING place="6" resultid="985" />
                    <RANKING place="2" resultid="986" />
                    <RANKING place="1" resultid="987" />
                    <RANKING place="4" resultid="988" />
                    <RANKING place="7" resultid="989" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6" agemax="11" agemin="11" name="Jahrgang 2012 - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="1" resultid="772" />
                    <RANKING place="3" resultid="773" />
                    <RANKING place="2" resultid="983" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7" agemax="12" agemin="12" name="Jahrgang 2011 - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="1" resultid="279" />
                    <RANKING place="4" resultid="280" />
                    <RANKING place="5" resultid="418" />
                    <RANKING place="3" resultid="774" />
                    <RANKING place="2" resultid="984" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8" agemax="13" agemin="13" name="Jahrgang 2010 - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="1" resultid="417" />
                    <RANKING place="2" resultid="982" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9" agemax="14" agemin="14" name="Jahrgang 2009 - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="1" resultid="768" />
                    <RANKING place="2" resultid="770" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10" agemax="15" agemin="15" name="Jahrgang 2008 - Süddeutsche Wertung" />
                <AGEGROUP agegroupid="11" agemax="16" agemin="16" name="Jahrgang 2007 - Süddeutsche Wertung" />
                <AGEGROUP agegroupid="12" agemax="17" agemin="17" name="Jahrgang 2006 - Süddeutsche Wertung" />
                <AGEGROUP agegroupid="13" agemax="21" agemin="18" name="Juniorinnen - Süddeutsche Wertung" />
                <AGEGROUP agegroupid="14" agemax="28" agemin="3" name="Offene Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="7" resultid="279" />
                    <RANKING place="11" resultid="280" />
                    <RANKING place="15" resultid="281" />
                    <RANKING place="23" resultid="416" />
                    <RANKING place="2" resultid="417" />
                    <RANKING place="12" resultid="418" />
                    <RANKING place="1" resultid="768" />
                    <RANKING place="6" resultid="770" />
                    <RANKING place="3" resultid="772" />
                    <RANKING place="9" resultid="773" />
                    <RANKING place="10" resultid="774" />
                    <RANKING place="21" resultid="775" />
                    <RANKING place="17" resultid="776" />
                    <RANKING place="5" resultid="982" />
                    <RANKING place="4" resultid="983" />
                    <RANKING place="8" resultid="984" />
                    <RANKING place="18" resultid="985" />
                    <RANKING place="14" resultid="986" />
                    <RANKING place="13" resultid="987" />
                    <RANKING place="16" resultid="988" />
                    <RANKING place="20" resultid="989" />
                    <RANKING place="25" resultid="990" />
                    <RANKING place="22" resultid="991" />
                    <RANKING place="19" resultid="992" />
                    <RANKING place="24" resultid="993" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="19" agemax="28" agemin="3" name="Offene internationale Wertung">
                  <RANKINGS>
                    <RANKING place="7" resultid="279" />
                    <RANKING place="11" resultid="280" />
                    <RANKING place="15" resultid="281" />
                    <RANKING place="23" resultid="416" />
                    <RANKING place="2" resultid="417" />
                    <RANKING place="12" resultid="418" />
                    <RANKING place="1" resultid="768" />
                    <RANKING place="6" resultid="770" />
                    <RANKING place="3" resultid="772" />
                    <RANKING place="9" resultid="773" />
                    <RANKING place="10" resultid="774" />
                    <RANKING place="21" resultid="775" />
                    <RANKING place="17" resultid="776" />
                    <RANKING place="5" resultid="982" />
                    <RANKING place="4" resultid="983" />
                    <RANKING place="8" resultid="984" />
                    <RANKING place="18" resultid="985" />
                    <RANKING place="14" resultid="986" />
                    <RANKING place="13" resultid="987" />
                    <RANKING place="16" resultid="988" />
                    <RANKING place="20" resultid="989" />
                    <RANKING place="25" resultid="990" />
                    <RANKING place="22" resultid="991" />
                    <RANKING place="19" resultid="992" />
                    <RANKING place="24" resultid="993" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15" agemax="44" agemin="29" name="Master A - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="1" resultid="147" />
                    <RANKING place="2" resultid="769" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="16" agemax="54" agemin="45" name="Master B - Süddeutsche Wertung" />
                <AGEGROUP agegroupid="17" agemax="-1" agemin="55" name="Master C - Süddeutsche Wertung" />
                <AGEGROUP agegroupid="18" agemax="-1" agemin="29" name="Offene internationale Wertung Master">
                  <RANKINGS>
                    <RANKING place="1" resultid="147" />
                    <RANKING place="2" resultid="769" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="4" number="4" gender="M" round="TIM">
              <SWIMSTYLE stroke="BIFIN" relaycount="1" distance="100" />
              <FEE value="500" currency="EUR" />
              <HEATS>
                <HEAT heatid="4001" number="1" />
                <HEAT heatid="4002" number="2" />
                <HEAT heatid="4003" number="3" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="4" agemax="9" agemin="3" name="Jahrgang 2014 und jünger - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="3" resultid="3" />
                    <RANKING place="1" resultid="285" />
                    <RANKING place="2" resultid="781" />
                    <RANKING place="4" resultid="997" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="10" agemin="10" name="Jahrgang 2013 - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="1" resultid="2" />
                    <RANKING place="2" resultid="996" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6" agemax="11" agemin="11" name="Jahrgang 2012 - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="3" resultid="1" />
                    <RANKING place="1" resultid="284" />
                    <RANKING place="2" resultid="780" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7" agemax="12" agemin="12" name="Jahrgang 2011 - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="3" resultid="782" />
                    <RANKING place="1" resultid="994" />
                    <RANKING place="2" resultid="995" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8" agemax="13" agemin="13" name="Jahrgang 2010 - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="1" resultid="779" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9" agemax="14" agemin="14" name="Jahrgang 2009 - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="1" resultid="778" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10" agemax="15" agemin="15" name="Jahrgang 2008 - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="1" resultid="283" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11" agemax="16" agemin="16" name="Jahrgang 2007 - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="1" resultid="419" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="12" agemax="17" agemin="17" name="Jahrgang 2006 - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="1" resultid="174" />
                    <RANKING place="2" resultid="420" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="13" agemax="21" agemin="18" name="Junioren - Süddeutsche Wertung" />
                <AGEGROUP agegroupid="14" agemax="30" agemin="3" name="Offene Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="16" resultid="1" />
                    <RANKING place="14" resultid="2" />
                    <RANKING place="15" resultid="3" />
                    <RANKING place="2" resultid="174" />
                    <RANKING place="1" resultid="282" />
                    <RANKING place="5" resultid="283" />
                    <RANKING place="7" resultid="284" />
                    <RANKING place="11" resultid="285" />
                    <RANKING place="4" resultid="419" />
                    <RANKING place="3" resultid="420" />
                    <RANKING place="6" resultid="778" />
                    <RANKING place="8" resultid="779" />
                    <RANKING place="13" resultid="780" />
                    <RANKING place="12" resultid="781" />
                    <RANKING place="17" resultid="782" />
                    <RANKING place="9" resultid="994" />
                    <RANKING place="10" resultid="995" />
                    <RANKING place="18" resultid="996" />
                    <RANKING place="19" resultid="997" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="19" agemax="30" agemin="3" name="Offene internationale Wertung">
                  <RANKINGS>
                    <RANKING place="16" resultid="1" />
                    <RANKING place="14" resultid="2" />
                    <RANKING place="15" resultid="3" />
                    <RANKING place="2" resultid="174" />
                    <RANKING place="1" resultid="282" />
                    <RANKING place="5" resultid="283" />
                    <RANKING place="7" resultid="284" />
                    <RANKING place="11" resultid="285" />
                    <RANKING place="4" resultid="419" />
                    <RANKING place="3" resultid="420" />
                    <RANKING place="6" resultid="778" />
                    <RANKING place="8" resultid="779" />
                    <RANKING place="13" resultid="780" />
                    <RANKING place="12" resultid="781" />
                    <RANKING place="17" resultid="782" />
                    <RANKING place="9" resultid="994" />
                    <RANKING place="10" resultid="995" />
                    <RANKING place="18" resultid="996" />
                    <RANKING place="19" resultid="997" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15" agemax="44" agemin="29" name="Master A - Süddeutsche Wertung" />
                <AGEGROUP agegroupid="16" agemax="54" agemin="45" name="Master B - Süddeutsche Wertung" />
                <AGEGROUP agegroupid="17" agemax="-1" agemin="55" name="Master C - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="1" resultid="117" />
                    <RANKING place="2" resultid="421" />
                    <RANKING place="3" resultid="422" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="18" agemax="-1" agemin="29" name="Offene internationale Wertung Master">
                  <RANKINGS>
                    <RANKING place="2" resultid="117" />
                    <RANKING place="3" resultid="421" />
                    <RANKING place="4" resultid="422" />
                    <RANKING place="1" resultid="952" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="5" number="5" gender="F" round="TIM">
              <SWIMSTYLE stroke="IMMERSION" technique="DIVE" relaycount="1" distance="400" />
              <FEE value="500" currency="EUR" />
              <HEATS>
                <HEAT heatid="5001" number="1" />
                <HEAT heatid="5002" number="2" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="4" agemax="9" agemin="12" name="Jahrgang 2014 und jünger - Süddeutsche Wertung" />
                <AGEGROUP agegroupid="5" agemax="10" agemin="12" name="Jahrgang 2013 - Süddeutsche Wertung" />
                <AGEGROUP agegroupid="6" agemax="11" agemin="12" name="Jahrgang 2012 - Süddeutsche Wertung" />
                <AGEGROUP agegroupid="7" agemax="12" agemin="12" name="Jahrgang 2011 - Süddeutsche Wertung" />
                <AGEGROUP agegroupid="8" agemax="13" agemin="13" name="Jahrgang 2010 - Süddeutsche Wertung" />
                <AGEGROUP agegroupid="9" agemax="14" agemin="14" name="Jahrgang 2009 - Süddeutsche Wertung" />
                <AGEGROUP agegroupid="10" agemax="15" agemin="15" name="Jahrgang 2008 - Süddeutsche Wertung" />
                <AGEGROUP agegroupid="11" agemax="16" agemin="16" name="Jahrgang 2007 - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="1" resultid="1048" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="12" agemax="17" agemin="17" name="Jahrgang 2006 - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="1" resultid="329" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="13" agemax="21" agemin="18" name="Juniorinnen - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="3" resultid="472" />
                    <RANKING place="1" resultid="1046" />
                    <RANKING place="2" resultid="1047" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="14" agemax="28" agemin="12" name="Offene Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="1" resultid="162" />
                    <RANKING place="2" resultid="163" />
                    <RANKING place="7" resultid="329" />
                    <RANKING place="9" resultid="472" />
                    <RANKING place="8" resultid="685" />
                    <RANKING place="6" resultid="977" />
                    <RANKING place="3" resultid="1046" />
                    <RANKING place="4" resultid="1047" />
                    <RANKING place="5" resultid="1048" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="19" agemax="28" agemin="12" name="Offene internationale Wertung">
                  <RANKINGS>
                    <RANKING place="1" resultid="162" />
                    <RANKING place="2" resultid="163" />
                    <RANKING place="7" resultid="329" />
                    <RANKING place="9" resultid="472" />
                    <RANKING place="8" resultid="685" />
                    <RANKING place="6" resultid="977" />
                    <RANKING place="3" resultid="1046" />
                    <RANKING place="4" resultid="1047" />
                    <RANKING place="5" resultid="1048" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15" agemax="44" agemin="29" name="Master A - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="1" resultid="164" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="16" agemax="54" agemin="45" name="Master B - Süddeutsche Wertung" />
                <AGEGROUP agegroupid="17" agemax="-1" agemin="55" name="Master C - Süddeutsche Wertung" />
                <AGEGROUP agegroupid="18" agemax="-1" agemin="29" name="Offene internationale Wertung Master">
                  <RANKINGS>
                    <RANKING place="1" resultid="164" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="6" number="6" gender="M" round="TIM">
              <SWIMSTYLE stroke="IMMERSION" technique="DIVE" relaycount="1" distance="400" />
              <FEE value="500" currency="EUR" />
              <HEATS>
                <HEAT heatid="6001" number="1" />
                <HEAT heatid="6002" number="2" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="4" agemax="9" agemin="12" name="Jahrgang 2014 und jünger - Süddeutsche Wertung" />
                <AGEGROUP agegroupid="5" agemax="10" agemin="12" name="Jahrgang 2013 - Süddeutsche Wertung" />
                <AGEGROUP agegroupid="6" agemax="11" agemin="12" name="Jahrgang 2012 - Süddeutsche Wertung" />
                <AGEGROUP agegroupid="7" agemax="12" agemin="12" name="Jahrgang 2011 - Süddeutsche Wertung" />
                <AGEGROUP agegroupid="8" agemax="13" agemin="13" name="Jahrgang 2010 - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="1" resultid="474" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9" agemax="14" agemin="14" name="Jahrgang 2009 - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="1" resultid="331" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10" agemax="15" agemin="15" name="Jahrgang 2008 - Süddeutsche Wertung" />
                <AGEGROUP agegroupid="11" agemax="16" agemin="16" name="Jahrgang 2007 - Süddeutsche Wertung" />
                <AGEGROUP agegroupid="12" agemax="17" agemin="17" name="Jahrgang 2006 - Süddeutsche Wertung" />
                <AGEGROUP agegroupid="13" agemax="21" agemin="18" name="Junioren - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="1" resultid="475" />
                    <RANKING place="2" resultid="686" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="14" agemax="28" agemin="12" name="Offene Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="3" resultid="331" />
                    <RANKING place="4" resultid="474" />
                    <RANKING place="1" resultid="475" />
                    <RANKING place="2" resultid="686" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="19" agemax="28" agemin="12" name="Offene internationale Wertung">
                  <RANKINGS>
                    <RANKING place="1" resultid="95" />
                    <RANKING place="5" resultid="331" />
                    <RANKING place="6" resultid="474" />
                    <RANKING place="2" resultid="475" />
                    <RANKING place="3" resultid="663" />
                    <RANKING place="4" resultid="686" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15" agemax="44" agemin="29" name="Master A - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="1" resultid="165" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="16" agemax="54" agemin="45" name="Master B - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="1" resultid="866" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="17" agemax="-1" agemin="55" name="Master C - Süddeutsche Wertung" />
                <AGEGROUP agegroupid="18" agemax="-1" agemin="29" name="Offene internationale Wertung Master">
                  <RANKINGS>
                    <RANKING place="1" resultid="165" />
                    <RANKING place="2" resultid="866" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="7" number="7" gender="F" round="TIM">
              <SWIMSTYLE stroke="APNEA" relaycount="1" distance="50" />
              <FEE value="500" currency="EUR" />
              <HEATS>
                <HEAT heatid="7001" number="1" />
                <HEAT heatid="7002" number="2" />
                <HEAT heatid="7003" number="3" />
                <HEAT heatid="7004" number="4" />
                <HEAT heatid="7005" number="5" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="4" agemax="9" agemin="14" name="Jahrgang 2014 und jünger - Süddeutsche Wertung" />
                <AGEGROUP agegroupid="5" agemax="10" agemin="14" name="Jahrgang 2013 - Süddeutsche Wertung" />
                <AGEGROUP agegroupid="6" agemax="11" agemin="14" name="Jahrgang 2012 - Süddeutsche Wertung" />
                <AGEGROUP agegroupid="7" agemax="12" agemin="14" name="Jahrgang 2011 - Süddeutsche Wertung" />
                <AGEGROUP agegroupid="8" agemax="13" agemin="14" name="Jahrgang 2010 - Süddeutsche Wertung" />
                <AGEGROUP agegroupid="9" agemax="14" agemin="14" name="Jahrgang 2009 - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="2" resultid="241" />
                    <RANKING place="6" resultid="245" />
                    <RANKING place="4" resultid="341" />
                    <RANKING place="5" resultid="689" />
                    <RANKING place="1" resultid="879" />
                    <RANKING place="3" resultid="884" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10" agemax="15" agemin="15" name="Jahrgang 2008 - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="1" resultid="242" />
                    <RANKING place="2" resultid="743" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11" agemax="16" agemin="16" name="Jahrgang 2007 - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="4" resultid="41" />
                    <RANKING place="3" resultid="69" />
                    <RANKING place="2" resultid="139" />
                    <RANKING place="1" resultid="1053" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="12" agemax="17" agemin="17" name="Jahrgang 2006 - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="1" resultid="339" />
                    <RANKING place="2" resultid="340" />
                    <RANKING place="5" resultid="688" />
                    <RANKING place="4" resultid="742" />
                    <RANKING place="3" resultid="881" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="13" agemax="21" agemin="18" name="Juniorinnen - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="1" resultid="138" />
                    <RANKING place="3" resultid="239" />
                    <RANKING place="6" resultid="240" />
                    <RANKING place="5" resultid="338" />
                    <RANKING place="8" resultid="483" />
                    <RANKING place="4" resultid="485" />
                    <RANKING place="9" resultid="882" />
                    <RANKING place="2" resultid="1052" />
                    <RANKING place="7" resultid="1054" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="14" agemax="28" agemin="14" name="Offene Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="29" resultid="41" />
                    <RANKING place="20" resultid="69" />
                    <RANKING place="1" resultid="138" />
                    <RANKING place="11" resultid="139" />
                    <RANKING place="8" resultid="166" />
                    <RANKING place="3" resultid="239" />
                    <RANKING place="9" resultid="240" />
                    <RANKING place="15" resultid="241" />
                    <RANKING place="13" resultid="242" />
                    <RANKING place="14" resultid="244" />
                    <RANKING place="27" resultid="245" />
                    <RANKING place="7" resultid="338" />
                    <RANKING place="16" resultid="339" />
                    <RANKING place="17" resultid="340" />
                    <RANKING place="24" resultid="341" />
                    <RANKING place="19" resultid="483" />
                    <RANKING place="4" resultid="485" />
                    <RANKING place="22" resultid="688" />
                    <RANKING place="26" resultid="689" />
                    <RANKING place="5" resultid="741" />
                    <RANKING place="21" resultid="742" />
                    <RANKING place="25" resultid="743" />
                    <RANKING place="10" resultid="879" />
                    <RANKING place="18" resultid="881" />
                    <RANKING place="28" resultid="882" />
                    <RANKING place="23" resultid="884" />
                    <RANKING place="2" resultid="1052" />
                    <RANKING place="6" resultid="1053" />
                    <RANKING place="12" resultid="1054" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="19" agemax="28" agemin="14" name="Offene internationale Wertung">
                  <RANKINGS>
                    <RANKING place="32" resultid="41" />
                    <RANKING place="22" resultid="69" />
                    <RANKING place="13" resultid="99" />
                    <RANKING place="1" resultid="138" />
                    <RANKING place="11" resultid="139" />
                    <RANKING place="8" resultid="166" />
                    <RANKING place="3" resultid="239" />
                    <RANKING place="9" resultid="240" />
                    <RANKING place="16" resultid="241" />
                    <RANKING place="14" resultid="242" />
                    <RANKING place="15" resultid="244" />
                    <RANKING place="30" resultid="245" />
                    <RANKING place="7" resultid="338" />
                    <RANKING place="17" resultid="339" />
                    <RANKING place="19" resultid="340" />
                    <RANKING place="26" resultid="341" />
                    <RANKING place="18" resultid="404" />
                    <RANKING place="28" resultid="405" />
                    <RANKING place="21" resultid="483" />
                    <RANKING place="4" resultid="485" />
                    <RANKING place="24" resultid="688" />
                    <RANKING place="29" resultid="689" />
                    <RANKING place="5" resultid="741" />
                    <RANKING place="23" resultid="742" />
                    <RANKING place="27" resultid="743" />
                    <RANKING place="10" resultid="879" />
                    <RANKING place="20" resultid="881" />
                    <RANKING place="31" resultid="882" />
                    <RANKING place="25" resultid="884" />
                    <RANKING place="2" resultid="1052" />
                    <RANKING place="6" resultid="1053" />
                    <RANKING place="12" resultid="1054" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15" agemax="44" agemin="29" name="Master A - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="1" resultid="883" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="16" agemax="54" agemin="45" name="Master B - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="1" resultid="486" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="17" agemax="-1" agemin="55" name="Master C - Süddeutsche Wertung" />
                <AGEGROUP agegroupid="18" agemax="-1" agemin="29" name="Offene internationale Wertung Master">
                  <RANKINGS>
                    <RANKING place="1" resultid="486" />
                    <RANKING place="2" resultid="883" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="8" number="8" gender="M" round="TIM">
              <SWIMSTYLE stroke="APNEA" relaycount="1" distance="50" />
              <FEE value="500" currency="EUR" />
              <HEATS>
                <HEAT heatid="8001" number="1" />
                <HEAT heatid="8002" number="2" />
                <HEAT heatid="8003" number="3" />
                <HEAT heatid="8004" number="4" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="4" agemax="9" agemin="14" name="Jahrgang 2014 und jünger - Süddeutsche Wertung" />
                <AGEGROUP agegroupid="5" agemax="10" agemin="14" name="Jahrgang 2013 - Süddeutsche Wertung" />
                <AGEGROUP agegroupid="6" agemax="11" agemin="14" name="Jahrgang 2012 - Süddeutsche Wertung" />
                <AGEGROUP agegroupid="7" agemax="12" agemin="14" name="Jahrgang 2011 - Süddeutsche Wertung" />
                <AGEGROUP agegroupid="8" agemax="13" agemin="14" name="Jahrgang 2010 - Süddeutsche Wertung" />
                <AGEGROUP agegroupid="9" agemax="14" agemin="14" name="Jahrgang 2009 - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="2" resultid="42" />
                    <RANKING place="3" resultid="44" />
                    <RANKING place="1" resultid="345" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10" agemax="15" agemin="15" name="Jahrgang 2008 - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="1" resultid="887" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11" agemax="16" agemin="16" name="Jahrgang 2007 - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="1" resultid="745" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="12" agemax="17" agemin="17" name="Jahrgang 2006 - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="4" resultid="43" />
                    <RANKING place="2" resultid="248" />
                    <RANKING place="3" resultid="490" />
                    <RANKING place="1" resultid="885" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="13" agemax="21" agemin="18" name="Junioren - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="2" resultid="246" />
                    <RANKING place="5" resultid="249" />
                    <RANKING place="3" resultid="487" />
                    <RANKING place="1" resultid="488" />
                    <RANKING place="4" resultid="491" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="14" agemax="28" agemin="14" name="Offene Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="15" resultid="42" />
                    <RANKING place="11" resultid="43" />
                    <RANKING place="16" resultid="44" />
                    <RANKING place="5" resultid="246" />
                    <RANKING place="7" resultid="248" />
                    <RANKING place="10" resultid="249" />
                    <RANKING place="4" resultid="342" />
                    <RANKING place="13" resultid="345" />
                    <RANKING place="6" resultid="487" />
                    <RANKING place="3" resultid="488" />
                    <RANKING place="8" resultid="490" />
                    <RANKING place="9" resultid="491" />
                    <RANKING place="2" resultid="744" />
                    <RANKING place="12" resultid="745" />
                    <RANKING place="1" resultid="885" />
                    <RANKING place="14" resultid="887" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="19" agemax="28" agemin="14" name="Offene internationale Wertung">
                  <RANKINGS>
                    <RANKING place="19" resultid="42" />
                    <RANKING place="15" resultid="43" />
                    <RANKING place="21" resultid="44" />
                    <RANKING place="9" resultid="101" />
                    <RANKING place="10" resultid="102" />
                    <RANKING place="6" resultid="246" />
                    <RANKING place="11" resultid="248" />
                    <RANKING place="14" resultid="249" />
                    <RANKING place="5" resultid="342" />
                    <RANKING place="17" resultid="345" />
                    <RANKING place="7" resultid="406" />
                    <RANKING place="20" resultid="407" />
                    <RANKING place="8" resultid="487" />
                    <RANKING place="4" resultid="488" />
                    <RANKING place="12" resultid="490" />
                    <RANKING place="13" resultid="491" />
                    <RANKING place="1" resultid="664" />
                    <RANKING place="3" resultid="744" />
                    <RANKING place="16" resultid="745" />
                    <RANKING place="2" resultid="885" />
                    <RANKING place="18" resultid="887" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15" agemax="44" agemin="29" name="Master A - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="1" resultid="167" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="16" agemax="54" agemin="45" name="Master B - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="1" resultid="344" />
                    <RANKING place="2" resultid="886" />
                    <RANKING place="4" resultid="888" />
                    <RANKING place="3" resultid="965" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="17" agemax="-1" agemin="55" name="Master C - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="2" resultid="119" />
                    <RANKING place="1" resultid="493" />
                    <RANKING place="3" resultid="494" />
                    <RANKING place="4" resultid="495" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="18" agemax="-1" agemin="29" name="Offene internationale Wertung Master">
                  <RANKINGS>
                    <RANKING place="7" resultid="119" />
                    <RANKING place="1" resultid="167" />
                    <RANKING place="2" resultid="344" />
                    <RANKING place="4" resultid="493" />
                    <RANKING place="8" resultid="494" />
                    <RANKING place="9" resultid="495" />
                    <RANKING place="3" resultid="886" />
                    <RANKING place="6" resultid="888" />
                    <RANKING place="5" resultid="965" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="9" number="9" gender="F" round="TIM">
              <SWIMSTYLE stroke="IMMERSION" technique="DIVE" relaycount="1" distance="50" />
              <FEE value="500" currency="EUR" />
              <HEATS>
                <HEAT heatid="9001" number="1" />
                <HEAT heatid="9002" number="2" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="4" agemax="9" agemin="12" name="Jahrgang 2014 und jünger - Süddeutsche Wertung" />
                <AGEGROUP agegroupid="5" agemax="10" agemin="12" name="Jahrgang 2013 - Süddeutsche Wertung" />
                <AGEGROUP agegroupid="6" agemax="11" agemin="12" name="Jahrgang 2012 - Süddeutsche Wertung" />
                <AGEGROUP agegroupid="7" agemax="12" agemin="12" name="Jahrgang 2011 - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="2" resultid="375" />
                    <RANKING place="1" resultid="944" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8" agemax="13" agemin="13" name="Jahrgang 2010 - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="3" resultid="762" />
                    <RANKING place="4" resultid="763" />
                    <RANKING place="1" resultid="945" />
                    <RANKING place="2" resultid="1096" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9" agemax="13" agemin="14" name="Jahrgang 2009 - Süddeutsche Wertung" />
                <AGEGROUP agegroupid="10" agemax="13" agemin="15" name="Jahrgang 2008 - Süddeutsche Wertung" />
                <AGEGROUP agegroupid="11" agemax="13" agemin="16" name="Jahrgang 2007 - Süddeutsche Wertung" />
                <AGEGROUP agegroupid="12" agemax="13" agemin="17" name="Jahrgang 2006 - Süddeutsche Wertung" />
                <AGEGROUP agegroupid="13" agemax="13" agemin="18" name="Juniorinnen - Süddeutsche Wertung" />
                <AGEGROUP agegroupid="14" agemax="13" agemin="12" name="Offene Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="6" resultid="375" />
                    <RANKING place="3" resultid="762" />
                    <RANKING place="5" resultid="763" />
                    <RANKING place="4" resultid="944" />
                    <RANKING place="1" resultid="945" />
                    <RANKING place="2" resultid="1096" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="19" agemax="13" agemin="12" name="Offene internationale Wertung">
                  <RANKINGS>
                    <RANKING place="8" resultid="375" />
                    <RANKING place="2" resultid="414" />
                    <RANKING place="4" resultid="415" />
                    <RANKING place="5" resultid="762" />
                    <RANKING place="7" resultid="763" />
                    <RANKING place="6" resultid="944" />
                    <RANKING place="1" resultid="945" />
                    <RANKING place="3" resultid="1096" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15" agemax="13" agemin="29" name="Master A - Süddeutsche Wertung" />
                <AGEGROUP agegroupid="16" agemax="13" agemin="45" name="Master B - Süddeutsche Wertung" />
                <AGEGROUP agegroupid="17" agemax="13" agemin="55" name="Master C - Süddeutsche Wertung" />
                <AGEGROUP agegroupid="18" agemax="13" agemin="29" name="Offene internationale Wertung Master" />
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="10" number="10" gender="M" round="TIM">
              <SWIMSTYLE stroke="IMMERSION" technique="DIVE" relaycount="1" distance="50" />
              <FEE value="500" currency="EUR" />
              <HEATS>
                <HEAT heatid="10001" number="1" />
                <HEAT heatid="10002" number="2" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="4" agemax="9" agemin="12" name="Jahrgang 2014 und jünger - Süddeutsche Wertung" />
                <AGEGROUP agegroupid="5" agemax="10" agemin="12" name="Jahrgang 2013 - Süddeutsche Wertung" />
                <AGEGROUP agegroupid="6" agemax="11" agemin="12" name="Jahrgang 2012 - Süddeutsche Wertung" />
                <AGEGROUP agegroupid="7" agemax="12" agemin="12" name="Jahrgang 2011 - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="1" resultid="277" />
                    <RANKING place="3" resultid="376" />
                    <RANKING place="2" resultid="537" />
                    <RANKING place="4" resultid="764" />
                    <RANKING place="6" resultid="1097" />
                    <RANKING place="5" resultid="1098" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8" agemax="13" agemin="13" name="Jahrgang 2010 - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="1" resultid="536" />
                    <RANKING place="2" resultid="948" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9" agemax="13" agemin="14" name="Jahrgang 2009 - Süddeutsche Wertung" />
                <AGEGROUP agegroupid="10" agemax="13" agemin="15" name="Jahrgang 2008 - Süddeutsche Wertung" />
                <AGEGROUP agegroupid="11" agemax="13" agemin="16" name="Jahrgang 2007 - Süddeutsche Wertung" />
                <AGEGROUP agegroupid="12" agemax="13" agemin="17" name="Jahrgang 2006 - Süddeutsche Wertung" />
                <AGEGROUP agegroupid="13" agemax="13" agemin="18" name="Junioren - Süddeutsche Wertung" />
                <AGEGROUP agegroupid="14" agemax="13" agemin="12" name="Offene Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="1" resultid="277" />
                    <RANKING place="5" resultid="376" />
                    <RANKING place="2" resultid="536" />
                    <RANKING place="3" resultid="537" />
                    <RANKING place="6" resultid="764" />
                    <RANKING place="4" resultid="948" />
                    <RANKING place="8" resultid="1097" />
                    <RANKING place="7" resultid="1098" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="19" agemax="13" agemin="12" name="Offene internationale Wertung">
                  <RANKINGS>
                    <RANKING place="1" resultid="277" />
                    <RANKING place="5" resultid="376" />
                    <RANKING place="2" resultid="536" />
                    <RANKING place="3" resultid="537" />
                    <RANKING place="6" resultid="764" />
                    <RANKING place="4" resultid="948" />
                    <RANKING place="8" resultid="1097" />
                    <RANKING place="7" resultid="1098" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15" agemax="13" agemin="29" name="Master A - Süddeutsche Wertung" />
                <AGEGROUP agegroupid="16" agemax="13" agemin="45" name="Master B - Süddeutsche Wertung" />
                <AGEGROUP agegroupid="17" agemax="13" agemin="55" name="Master C - Süddeutsche Wertung" />
                <AGEGROUP agegroupid="18" agemax="13" agemin="29" name="Offene internationale Wertung Master" />
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="11" number="11" gender="F" round="TIM">
              <SWIMSTYLE stroke="SURFACE" relaycount="1" distance="200" />
              <FEE value="500" currency="EUR" />
              <HEATS>
                <HEAT heatid="11001" number="1" />
                <HEAT heatid="11002" number="2" />
                <HEAT heatid="11003" number="3" />
                <HEAT heatid="11004" number="4" />
                <HEAT heatid="11005" number="5" />
                <HEAT heatid="11006" number="6" />
                <HEAT heatid="11007" number="7" />
                <HEAT heatid="11008" number="8" />
                <HEAT heatid="11009" number="9" />
                <HEAT heatid="11010" number="10" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="4" agemax="9" agemin="3" name="Jahrgang 2014 und jünger - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="4" resultid="210" />
                    <RANKING place="1" resultid="313" />
                    <RANKING place="2" resultid="463" />
                    <RANKING place="3" resultid="1021" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="10" agemin="10" name="Jahrgang 2013 - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="5" resultid="311" />
                    <RANKING place="7" resultid="461" />
                    <RANKING place="10" resultid="833" />
                    <RANKING place="9" resultid="834" />
                    <RANKING place="1" resultid="1026" />
                    <RANKING place="4" resultid="1027" />
                    <RANKING place="3" resultid="1028" />
                    <RANKING place="2" resultid="1029" />
                    <RANKING place="6" resultid="1030" />
                    <RANKING place="8" resultid="1031" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6" agemax="11" agemin="11" name="Jahrgang 2012 - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="2" resultid="207" />
                    <RANKING place="3" resultid="208" />
                    <RANKING place="9" resultid="456" />
                    <RANKING place="6" resultid="724" />
                    <RANKING place="4" resultid="828" />
                    <RANKING place="5" resultid="829" />
                    <RANKING place="8" resultid="830" />
                    <RANKING place="7" resultid="832" />
                    <RANKING place="1" resultid="1023" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7" agemax="12" agemin="12" name="Jahrgang 2011 - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="1" resultid="133" />
                    <RANKING place="5" resultid="209" />
                    <RANKING place="4" resultid="309" />
                    <RANKING place="7" resultid="310" />
                    <RANKING place="10" resultid="312" />
                    <RANKING place="9" resultid="460" />
                    <RANKING place="8" resultid="726" />
                    <RANKING place="2" resultid="827" />
                    <RANKING place="6" resultid="831" />
                    <RANKING place="3" resultid="1025" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8" agemax="13" agemin="13" name="Jahrgang 2010 - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="3" resultid="134" />
                    <RANKING place="2" resultid="458" />
                    <RANKING place="6" resultid="459" />
                    <RANKING place="4" resultid="723" />
                    <RANKING place="7" resultid="725" />
                    <RANKING place="8" resultid="819" />
                    <RANKING place="1" resultid="822" />
                    <RANKING place="5" resultid="1024" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9" agemax="14" agemin="14" name="Jahrgang 2009 - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="7" resultid="66" />
                    <RANKING place="2" resultid="205" />
                    <RANKING place="5" resultid="206" />
                    <RANKING place="4" resultid="676" />
                    <RANKING place="1" resultid="820" />
                    <RANKING place="3" resultid="823" />
                    <RANKING place="6" resultid="826" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10" agemax="15" agemin="15" name="Jahrgang 2008 - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="1" resultid="721" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11" agemax="16" agemin="16" name="Jahrgang 2007 - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="2" resultid="135" />
                    <RANKING place="1" resultid="1022" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="12" agemax="17" agemin="17" name="Jahrgang 2006 - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="1" resultid="307" />
                    <RANKING place="3" resultid="677" />
                    <RANKING place="2" resultid="821" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="13" agemax="21" agemin="18" name="Juniorinnen - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="1" resultid="132" />
                    <RANKING place="3" resultid="204" />
                    <RANKING place="2" resultid="306" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="14" agemax="28" agemin="3" name="Offene Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="11" resultid="20" />
                    <RANKING place="39" resultid="66" />
                    <RANKING place="1" resultid="132" />
                    <RANKING place="26" resultid="133" />
                    <RANKING place="20" resultid="134" />
                    <RANKING place="33" resultid="135" />
                    <RANKING place="2" resultid="155" />
                    <RANKING place="4" resultid="204" />
                    <RANKING place="7" resultid="205" />
                    <RANKING place="18" resultid="206" />
                    <RANKING place="22" resultid="207" />
                    <RANKING place="24" resultid="208" />
                    <RANKING place="30" resultid="209" />
                    <RANKING place="60" resultid="210" />
                    <RANKING place="3" resultid="306" />
                    <RANKING place="10" resultid="307" />
                    <RANKING place="29" resultid="309" />
                    <RANKING place="41" resultid="310" />
                    <RANKING place="50" resultid="311" />
                    <RANKING place="52" resultid="312" />
                    <RANKING place="54" resultid="313" />
                    <RANKING place="44" resultid="456" />
                    <RANKING place="16" resultid="458" />
                    <RANKING place="31" resultid="459" />
                    <RANKING place="47" resultid="460" />
                    <RANKING place="53" resultid="461" />
                    <RANKING place="55" resultid="463" />
                    <RANKING place="8" resultid="675" />
                    <RANKING place="17" resultid="676" />
                    <RANKING place="15" resultid="677" />
                    <RANKING place="13" resultid="721" />
                    <RANKING place="23" resultid="723" />
                    <RANKING place="36" resultid="724" />
                    <RANKING place="35" resultid="725" />
                    <RANKING place="45" resultid="726" />
                    <RANKING place="46" resultid="819" />
                    <RANKING place="6" resultid="820" />
                    <RANKING place="12" resultid="821" />
                    <RANKING place="9" resultid="822" />
                    <RANKING place="14" resultid="823" />
                    <RANKING place="21" resultid="826" />
                    <RANKING place="27" resultid="827" />
                    <RANKING place="32" resultid="828" />
                    <RANKING place="34" resultid="829" />
                    <RANKING place="42" resultid="830" />
                    <RANKING place="37" resultid="831" />
                    <RANKING place="38" resultid="832" />
                    <RANKING place="59" resultid="833" />
                    <RANKING place="58" resultid="834" />
                    <RANKING place="56" resultid="1021" />
                    <RANKING place="5" resultid="1022" />
                    <RANKING place="19" resultid="1023" />
                    <RANKING place="25" resultid="1024" />
                    <RANKING place="28" resultid="1025" />
                    <RANKING place="40" resultid="1026" />
                    <RANKING place="49" resultid="1027" />
                    <RANKING place="48" resultid="1028" />
                    <RANKING place="43" resultid="1029" />
                    <RANKING place="51" resultid="1030" />
                    <RANKING place="57" resultid="1031" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="19" agemax="28" agemin="3" name="Offene internationale Wertung">
                  <RANKINGS>
                    <RANKING place="12" resultid="20" />
                    <RANKING place="47" resultid="66" />
                    <RANKING place="11" resultid="83" />
                    <RANKING place="22" resultid="84" />
                    <RANKING place="1" resultid="132" />
                    <RANKING place="33" resultid="133" />
                    <RANKING place="25" resultid="134" />
                    <RANKING place="41" resultid="135" />
                    <RANKING place="2" resultid="155" />
                    <RANKING place="4" resultid="204" />
                    <RANKING place="7" resultid="205" />
                    <RANKING place="23" resultid="206" />
                    <RANKING place="29" resultid="207" />
                    <RANKING place="31" resultid="208" />
                    <RANKING place="38" resultid="209" />
                    <RANKING place="68" resultid="210" />
                    <RANKING place="3" resultid="306" />
                    <RANKING place="10" resultid="307" />
                    <RANKING place="37" resultid="309" />
                    <RANKING place="49" resultid="310" />
                    <RANKING place="58" resultid="311" />
                    <RANKING place="60" resultid="312" />
                    <RANKING place="62" resultid="313" />
                    <RANKING place="14" resultid="392" />
                    <RANKING place="13" resultid="393" />
                    <RANKING place="27" resultid="394" />
                    <RANKING place="20" resultid="395" />
                    <RANKING place="52" resultid="456" />
                    <RANKING place="19" resultid="458" />
                    <RANKING place="39" resultid="459" />
                    <RANKING place="55" resultid="460" />
                    <RANKING place="61" resultid="461" />
                    <RANKING place="63" resultid="463" />
                    <RANKING place="28" resultid="659" />
                    <RANKING place="34" resultid="660" />
                    <RANKING place="8" resultid="675" />
                    <RANKING place="21" resultid="676" />
                    <RANKING place="18" resultid="677" />
                    <RANKING place="16" resultid="721" />
                    <RANKING place="30" resultid="723" />
                    <RANKING place="44" resultid="724" />
                    <RANKING place="43" resultid="725" />
                    <RANKING place="53" resultid="726" />
                    <RANKING place="54" resultid="819" />
                    <RANKING place="6" resultid="820" />
                    <RANKING place="15" resultid="821" />
                    <RANKING place="9" resultid="822" />
                    <RANKING place="17" resultid="823" />
                    <RANKING place="26" resultid="826" />
                    <RANKING place="35" resultid="827" />
                    <RANKING place="40" resultid="828" />
                    <RANKING place="42" resultid="829" />
                    <RANKING place="50" resultid="830" />
                    <RANKING place="45" resultid="831" />
                    <RANKING place="46" resultid="832" />
                    <RANKING place="67" resultid="833" />
                    <RANKING place="66" resultid="834" />
                    <RANKING place="64" resultid="1021" />
                    <RANKING place="5" resultid="1022" />
                    <RANKING place="24" resultid="1023" />
                    <RANKING place="32" resultid="1024" />
                    <RANKING place="36" resultid="1025" />
                    <RANKING place="48" resultid="1026" />
                    <RANKING place="57" resultid="1027" />
                    <RANKING place="56" resultid="1028" />
                    <RANKING place="51" resultid="1029" />
                    <RANKING place="59" resultid="1030" />
                    <RANKING place="65" resultid="1031" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15" agemax="44" agemin="29" name="Master A - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="3" resultid="156" />
                    <RANKING place="1" resultid="824" />
                    <RANKING place="2" resultid="959" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="16" agemax="54" agemin="45" name="Master B - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="1" resultid="457" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="17" agemax="-1" agemin="55" name="Master C - Süddeutsche Wertung" />
                <AGEGROUP agegroupid="18" agemax="-1" agemin="29" name="Offene internationale Wertung Master">
                  <RANKINGS>
                    <RANKING place="4" resultid="156" />
                    <RANKING place="1" resultid="457" />
                    <RANKING place="2" resultid="824" />
                    <RANKING place="3" resultid="959" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="12" number="12" gender="M" round="TIM">
              <SWIMSTYLE stroke="SURFACE" relaycount="1" distance="200" />
              <FEE value="500" currency="EUR" />
              <HEATS>
                <HEAT heatid="12001" number="1" />
                <HEAT heatid="12002" number="2" />
                <HEAT heatid="12003" number="3" />
                <HEAT heatid="12004" number="4" />
                <HEAT heatid="12005" number="5" />
                <HEAT heatid="12006" number="6" />
                <HEAT heatid="12007" number="7" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="4" agemax="9" agemin="3" name="Jahrgang 2014 und jünger - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="3" resultid="28" />
                    <RANKING place="1" resultid="320" />
                    <RANKING place="4" resultid="467" />
                    <RANKING place="2" resultid="844" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="10" agemin="10" name="Jahrgang 2013 - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="3" resultid="26" />
                    <RANKING place="1" resultid="214" />
                    <RANKING place="2" resultid="215" />
                    <RANKING place="4" resultid="1034" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6" agemax="11" agemin="11" name="Jahrgang 2012 - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="3" resultid="27" />
                    <RANKING place="1" resultid="213" />
                    <RANKING place="2" resultid="319" />
                    <RANKING place="4" resultid="681" />
                    <RANKING place="5" resultid="845" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7" agemax="12" agemin="12" name="Jahrgang 2011 - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="2" resultid="318" />
                    <RANKING place="1" resultid="466" />
                    <RANKING place="5" resultid="729" />
                    <RANKING place="6" resultid="730" />
                    <RANKING place="4" resultid="1032" />
                    <RANKING place="3" resultid="1033" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8" agemax="13" agemin="13" name="Jahrgang 2010 - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="1" resultid="837" />
                    <RANKING place="2" resultid="840" />
                    <RANKING place="3" resultid="842" />
                    <RANKING place="4" resultid="843" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9" agemax="14" agemin="14" name="Jahrgang 2009 - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="2" resultid="24" />
                    <RANKING place="4" resultid="25" />
                    <RANKING place="1" resultid="315" />
                    <RANKING place="5" resultid="465" />
                    <RANKING place="3" resultid="839" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10" agemax="15" agemin="15" name="Jahrgang 2008 - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="2" resultid="22" />
                    <RANKING place="1" resultid="314" />
                    <RANKING place="4" resultid="317" />
                    <RANKING place="3" resultid="838" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11" agemax="16" agemin="16" name="Jahrgang 2007 - Süddeutsche Wertung" />
                <AGEGROUP agegroupid="12" agemax="17" agemin="17" name="Jahrgang 2006 - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="2" resultid="23" />
                    <RANKING place="1" resultid="836" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="13" agemax="21" agemin="18" name="Junioren - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="3" resultid="212" />
                    <RANKING place="1" resultid="464" />
                    <RANKING place="2" resultid="679" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="14" agemax="28" agemin="3" name="Offene Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="7" resultid="22" />
                    <RANKING place="6" resultid="23" />
                    <RANKING place="12" resultid="24" />
                    <RANKING place="15" resultid="25" />
                    <RANKING place="30" resultid="26" />
                    <RANKING place="24" resultid="27" />
                    <RANKING place="35" resultid="28" />
                    <RANKING place="8" resultid="212" />
                    <RANKING place="21" resultid="213" />
                    <RANKING place="25" resultid="214" />
                    <RANKING place="28" resultid="215" />
                    <RANKING place="4" resultid="314" />
                    <RANKING place="10" resultid="315" />
                    <RANKING place="16" resultid="317" />
                    <RANKING place="20" resultid="318" />
                    <RANKING place="22" resultid="319" />
                    <RANKING place="31" resultid="320" />
                    <RANKING place="3" resultid="464" />
                    <RANKING place="19" resultid="465" />
                    <RANKING place="14" resultid="466" />
                    <RANKING place="38" resultid="467" />
                    <RANKING place="5" resultid="679" />
                    <RANKING place="27" resultid="681" />
                    <RANKING place="2" resultid="727" />
                    <RANKING place="32" resultid="729" />
                    <RANKING place="37" resultid="730" />
                    <RANKING place="1" resultid="836" />
                    <RANKING place="11" resultid="837" />
                    <RANKING place="9" resultid="838" />
                    <RANKING place="13" resultid="839" />
                    <RANKING place="17" resultid="840" />
                    <RANKING place="18" resultid="842" />
                    <RANKING place="29" resultid="843" />
                    <RANKING place="33" resultid="844" />
                    <RANKING place="34" resultid="845" />
                    <RANKING place="26" resultid="1032" />
                    <RANKING place="23" resultid="1033" />
                    <RANKING place="36" resultid="1034" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="19" agemax="28" agemin="3" name="Offene internationale Wertung">
                  <RANKINGS>
                    <RANKING place="11" resultid="22" />
                    <RANKING place="10" resultid="23" />
                    <RANKING place="17" resultid="24" />
                    <RANKING place="20" resultid="25" />
                    <RANKING place="35" resultid="26" />
                    <RANKING place="29" resultid="27" />
                    <RANKING place="40" resultid="28" />
                    <RANKING place="1" resultid="85" />
                    <RANKING place="6" resultid="86" />
                    <RANKING place="9" resultid="87" />
                    <RANKING place="8" resultid="88" />
                    <RANKING place="12" resultid="212" />
                    <RANKING place="26" resultid="213" />
                    <RANKING place="30" resultid="214" />
                    <RANKING place="33" resultid="215" />
                    <RANKING place="5" resultid="314" />
                    <RANKING place="15" resultid="315" />
                    <RANKING place="21" resultid="317" />
                    <RANKING place="25" resultid="318" />
                    <RANKING place="27" resultid="319" />
                    <RANKING place="36" resultid="320" />
                    <RANKING place="14" resultid="396" />
                    <RANKING place="4" resultid="464" />
                    <RANKING place="24" resultid="465" />
                    <RANKING place="19" resultid="466" />
                    <RANKING place="43" resultid="467" />
                    <RANKING place="7" resultid="679" />
                    <RANKING place="32" resultid="681" />
                    <RANKING place="3" resultid="727" />
                    <RANKING place="37" resultid="729" />
                    <RANKING place="42" resultid="730" />
                    <RANKING place="2" resultid="836" />
                    <RANKING place="16" resultid="837" />
                    <RANKING place="13" resultid="838" />
                    <RANKING place="18" resultid="839" />
                    <RANKING place="22" resultid="840" />
                    <RANKING place="23" resultid="842" />
                    <RANKING place="34" resultid="843" />
                    <RANKING place="38" resultid="844" />
                    <RANKING place="39" resultid="845" />
                    <RANKING place="31" resultid="1032" />
                    <RANKING place="28" resultid="1033" />
                    <RANKING place="41" resultid="1034" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15" agemax="44" agemin="29" name="Master A - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="1" resultid="157" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="16" agemax="54" agemin="45" name="Master B - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="2" resultid="316" />
                    <RANKING place="1" resultid="966" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="17" agemax="-1" agemin="55" name="Master C - Süddeutsche Wertung" />
                <AGEGROUP agegroupid="18" agemax="-1" agemin="29" name="Offene internationale Wertung Master">
                  <RANKINGS>
                    <RANKING place="1" resultid="157" />
                    <RANKING place="4" resultid="316" />
                    <RANKING place="2" resultid="954" />
                    <RANKING place="3" resultid="966" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="13" number="13" gender="X" round="TIM">
              <SWIMSTYLE stroke="SURFACE" relaycount="4" distance="50" />
              <FEE value="800" currency="EUR" />
              <HEATS>
                <HEAT heatid="13001" number="1" />
                <HEAT heatid="13002" number="2" />
                <HEAT heatid="13003" number="3" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="2" agemax="11" agemin="3" name="Kategorie S3 - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="1" resultid="238" />
                    <RANKING place="3" resultid="876" />
                    <RANKING place="4" resultid="877" />
                    <RANKING place="2" resultid="1051" />
                    <RANKING place="5" resultid="1101" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3" agemax="14" agemin="12" name="Kategorie S2 - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="5" resultid="337" />
                    <RANKING place="2" resultid="481" />
                    <RANKING place="1" resultid="874" />
                    <RANKING place="3" resultid="875" />
                    <RANKING place="6" resultid="970" />
                    <RANKING place="4" resultid="1050" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="17" agemin="15" name="Kategorie S1 - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="1" resultid="237" />
                    <RANKING place="2" resultid="336" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7" agemax="28" agemin="3" name="Offene Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="8" resultid="40" />
                    <RANKING place="5" resultid="237" />
                    <RANKING place="11" resultid="238" />
                    <RANKING place="1" resultid="335" />
                    <RANKING place="7" resultid="336" />
                    <RANKING place="13" resultid="337" />
                    <RANKING place="2" resultid="480" />
                    <RANKING place="9" resultid="481" />
                    <RANKING place="4" resultid="873" />
                    <RANKING place="6" resultid="874" />
                    <RANKING place="10" resultid="875" />
                    <RANKING place="16" resultid="876" />
                    <RANKING place="17" resultid="877" />
                    <RANKING place="3" resultid="969" />
                    <RANKING place="14" resultid="970" />
                    <RANKING place="12" resultid="1050" />
                    <RANKING place="15" resultid="1051" />
                    <RANKING place="18" resultid="1101" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11" agemax="28" agemin="3" name="Offene internationale Wertung">
                  <RANKINGS>
                    <RANKING place="10" resultid="40" />
                    <RANKING place="3" resultid="98" />
                    <RANKING place="6" resultid="237" />
                    <RANKING place="13" resultid="238" />
                    <RANKING place="1" resultid="335" />
                    <RANKING place="9" resultid="336" />
                    <RANKING place="15" resultid="337" />
                    <RANKING place="7" resultid="403" />
                    <RANKING place="2" resultid="480" />
                    <RANKING place="11" resultid="481" />
                    <RANKING place="5" resultid="873" />
                    <RANKING place="8" resultid="874" />
                    <RANKING place="12" resultid="875" />
                    <RANKING place="18" resultid="876" />
                    <RANKING place="19" resultid="877" />
                    <RANKING place="4" resultid="969" />
                    <RANKING place="16" resultid="970" />
                    <RANKING place="14" resultid="1050" />
                    <RANKING place="17" resultid="1051" />
                    <RANKING place="20" resultid="1101" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8" agemax="28" agemin="176" easy.ak="176" calculate="TOTAL" name="Masters A - Süddeutsche Wertung" />
                <AGEGROUP agegroupid="9" agemax="28" agemin="400" easy.ak="400" calculate="TOTAL" name="Masters B - Süddeutsche Wertung" />
                <AGEGROUP agegroupid="10" agemax="28" agemin="400" easy.ak="400" calculate="TOTAL" name="Offene internationale Wertung Master" />
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="14" number="14" gender="X" round="TIM">
              <SWIMSTYLE stroke="SURFACE" relaycount="4" distance="50" />
              <FEE value="800" currency="EUR" />
              <HEATS>
                <HEAT heatid="14001" number="1" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="2" agemax="11" agemin="29" name="Kategorie S3 - Süddeutsche Wertung" />
                <AGEGROUP agegroupid="3" agemax="14" agemin="29" name="Kategorie S2 - Süddeutsche Wertung" />
                <AGEGROUP agegroupid="4" agemax="17" agemin="29" name="Kategorie S1 - Süddeutsche Wertung" />
                <AGEGROUP agegroupid="7" agemax="123" agemin="29" name="Offene Süddeutsche Wertung" />
                <AGEGROUP agegroupid="11" agemax="123" agemin="29" name="Offene internationale Wertung" />
                <AGEGROUP agegroupid="8" agemax="-1" agemin="176" easy.ak="176" calculate="TOTAL" name="Masters A - Süddeutsche Wertung" />
                <AGEGROUP agegroupid="9" agemax="-1" agemin="400" easy.ak="400" calculate="TOTAL" name="Masters B - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="2" resultid="482" />
                    <RANKING place="1" resultid="878" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10" agemax="-1" agemin="400" easy.ak="400" calculate="TOTAL" name="Offene internationale Wertung Master">
                  <RANKINGS>
                    <RANKING place="2" resultid="482" />
                    <RANKING place="1" resultid="878" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="15" number="15" gender="X" round="TIM">
              <SWIMSTYLE stroke="SURFACE" relaycount="1" distance="1500" />
              <FEE value="500" currency="EUR" />
              <HEATS>
                <HEAT heatid="15001" number="1" />
                <HEAT heatid="15002" number="2" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="4" agemax="9" agemin="12" name="weiblich: Jahrgang 2014 und jünger - Süddeutsche Wertung" />
                <AGEGROUP agegroupid="5" agemax="10" agemin="12" name="weiblich: Jahrgang 2013 - Süddeutsche Wertung" />
                <AGEGROUP agegroupid="6" agemax="11" agemin="12" name="weiblich: Jahrgang 2012 - Süddeutsche Wertung" />
                <AGEGROUP agegroupid="7" agemax="12" agemin="12" name="weiblich: Jahrgang 2011 - Süddeutsche Wertung" />
                <AGEGROUP agegroupid="8" agemax="13" agemin="13" name="weiblich: Jahrgang 2010 - Süddeutsche Wertung" />
                <AGEGROUP agegroupid="9" agemax="14" agemin="14" name="weiblich: Jahrgang 2009 - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="1" resultid="818" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10" agemax="15" agemin="15" name="weiblich: Jahrgang 2008 - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="1" resultid="720" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11" agemax="16" agemin="16" name="weiblich: Jahrgang 2007 - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="2" resultid="65" />
                    <RANKING place="1" resultid="131" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="12" agemax="17" agemin="17" name="weiblich: Jahrgang 2006 - Süddeutsche Wertung" />
                <AGEGROUP agegroupid="13" agemax="21" agemin="18" name="Juniorinnen - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="1" resultid="1020" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="14" agemax="28" agemin="12" name="weiblich: Offene Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="6" resultid="19" />
                    <RANKING place="4" resultid="65" />
                    <RANKING place="2" resultid="131" />
                    <RANKING place="1" resultid="154" />
                    <RANKING place="7" resultid="720" />
                    <RANKING place="5" resultid="818" />
                    <RANKING place="3" resultid="1020" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="19" agemax="28" agemin="12" name="weiblich: Offene internationale Wertung">
                  <RANKINGS>
                    <RANKING place="6" resultid="19" />
                    <RANKING place="4" resultid="65" />
                    <RANKING place="2" resultid="131" />
                    <RANKING place="1" resultid="154" />
                    <RANKING place="7" resultid="720" />
                    <RANKING place="5" resultid="818" />
                    <RANKING place="3" resultid="1020" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15" agemax="28" agemin="29" name="weiblich: Master A - Süddeutsche Wertung" />
                <AGEGROUP agegroupid="16" agemax="28" agemin="45" name="weiblich: Master B - Süddeutsche Wertung" />
                <AGEGROUP agegroupid="17" agemax="28" agemin="55" name="weiblich: Master C - Süddeutsche Wertung" />
                <AGEGROUP agegroupid="18" agemax="28" agemin="29" name="weiblich: Offene internationale Wertung Master" />
                <AGEGROUP agegroupid="23" agemax="9" agemin="12" name="männlich: Jahrgang 2014 und jünger - Süddeutsche Wertung" />
                <AGEGROUP agegroupid="24" agemax="10" agemin="12" name="männlich: Jahrgang 2013 - Süddeutsche Wertung" />
                <AGEGROUP agegroupid="25" agemax="11" agemin="12" name="männlich: Jahrgang 2012 - Süddeutsche Wertung" />
                <AGEGROUP agegroupid="26" agemax="12" agemin="12" name="männlich: Jahrgang 2011 - Süddeutsche Wertung" />
                <AGEGROUP agegroupid="27" agemax="13" agemin="13" name="männlich: Jahrgang 2010 - Süddeutsche Wertung" />
                <AGEGROUP agegroupid="28" agemax="14" agemin="14" name="männlich: Jahrgang 2009 - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="1" resultid="817" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="29" agemax="15" agemin="15" name="männlich: Jahrgang 2008 - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="1" resultid="17" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="30" agemax="16" agemin="16" name="männlich: Jahrgang 2007 - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="1" resultid="719" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="31" agemax="17" agemin="17" name="männlich: Jahrgang 2006 - Süddeutsche Wertung" />
                <AGEGROUP agegroupid="32" agemax="21" agemin="18" name="Junioren - Süddeutsche Wertung" />
                <AGEGROUP agegroupid="33" agemax="28" agemin="12" name="männlich: Offene Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="1" resultid="17" />
                    <RANKING place="2" resultid="719" />
                    <RANKING place="3" resultid="817" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="38" agemax="28" agemin="12" name="männlich: Offene internationale Wertung">
                  <RANKINGS>
                    <RANKING place="1" resultid="17" />
                    <RANKING place="2" resultid="719" />
                    <RANKING place="3" resultid="817" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="34" agemax="28" agemin="29" name="männlich: Master A - Süddeutsche Wertung" />
                <AGEGROUP agegroupid="35" agemax="28" agemin="45" name="männlich: Master B - Süddeutsche Wertung" />
                <AGEGROUP agegroupid="36" agemax="28" agemin="55" name="männlich: Master C - Süddeutsche Wertung" />
                <AGEGROUP agegroupid="37" agemax="28" agemin="29" name="männlich: Offene internationale Wertung Master" />
              </AGEGROUPS>
            </EVENT>
          </EVENTS>
        </SESSION>
        <SESSION number="2" date="2023-03-26" daytime="09:10" officialmeeting="08:40" warmupfrom="08:00">
          <EVENTS>
            <EVENT eventid="16" number="16" gender="F" round="TIM">
              <SWIMSTYLE stroke="SURFACE" relaycount="1" distance="50" />
              <FEE value="500" currency="EUR" />
              <HEATS>
                <HEAT heatid="16001" number="1" />
                <HEAT heatid="16002" number="2" />
                <HEAT heatid="16003" number="3" />
                <HEAT heatid="16004" number="4" />
                <HEAT heatid="16005" number="5" />
                <HEAT heatid="16006" number="6" />
                <HEAT heatid="16007" number="7" />
                <HEAT heatid="16008" number="8" />
                <HEAT heatid="16009" number="9" />
                <HEAT heatid="16010" number="10" />
                <HEAT heatid="16011" number="11" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="4" agemax="9" agemin="3" name="Jahrgang 2014 und jünger - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="1" resultid="268" />
                    <RANKING place="1" resultid="368" />
                    <RANKING place="3" resultid="525" />
                    <RANKING place="4" resultid="756" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="10" agemin="10" name="Jahrgang 2013 - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="6" resultid="367" />
                    <RANKING place="7" resultid="524" />
                    <RANKING place="1" resultid="1086" />
                    <RANKING place="2" resultid="1087" />
                    <RANKING place="3" resultid="1088" />
                    <RANKING place="5" resultid="1089" />
                    <RANKING place="4" resultid="1090" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6" agemax="11" agemin="11" name="Jahrgang 2012 - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="1" resultid="266" />
                    <RANKING place="8" resultid="522" />
                    <RANKING place="4" resultid="754" />
                    <RANKING place="5" resultid="927" />
                    <RANKING place="7" resultid="928" />
                    <RANKING place="6" resultid="931" />
                    <RANKING place="2" resultid="932" />
                    <RANKING place="3" resultid="1084" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7" agemax="12" agemin="12" name="Jahrgang 2011 - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="1" resultid="143" />
                    <RANKING place="4" resultid="267" />
                    <RANKING place="7" resultid="364" />
                    <RANKING place="6" resultid="365" />
                    <RANKING place="8" resultid="366" />
                    <RANKING place="2" resultid="519" />
                    <RANKING place="9" resultid="755" />
                    <RANKING place="3" resultid="924" />
                    <RANKING place="10" resultid="929" />
                    <RANKING place="5" resultid="1085" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8" agemax="13" agemin="13" name="Jahrgang 2010 - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="2" resultid="142" />
                    <RANKING place="4" resultid="518" />
                    <RANKING place="6" resultid="520" />
                    <RANKING place="5" resultid="752" />
                    <RANKING place="7" resultid="753" />
                    <RANKING place="1" resultid="918" />
                    <RANKING place="8" resultid="930" />
                    <RANKING place="3" resultid="1083" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9" agemax="14" agemin="14" name="Jahrgang 2009 - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="9" resultid="71" />
                    <RANKING place="3" resultid="260" />
                    <RANKING place="5" resultid="264" />
                    <RANKING place="6" resultid="363" />
                    <RANKING place="8" resultid="693" />
                    <RANKING place="1" resultid="915" />
                    <RANKING place="2" resultid="919" />
                    <RANKING place="4" resultid="921" />
                    <RANKING place="7" resultid="923" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10" agemax="15" agemin="15" name="Jahrgang 2008 - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="1" resultid="261" />
                    <RANKING place="2" resultid="749" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11" agemax="16" agemin="16" name="Jahrgang 2007 - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="4" resultid="50" />
                    <RANKING place="3" resultid="144" />
                    <RANKING place="2" resultid="926" />
                    <RANKING place="1" resultid="1082" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="12" agemax="17" agemin="17" name="Jahrgang 2006 - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="1" resultid="361" />
                    <RANKING place="2" resultid="362" />
                    <RANKING place="5" resultid="692" />
                    <RANKING place="4" resultid="750" />
                    <RANKING place="3" resultid="917" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="13" agemax="21" agemin="18" name="Juniorinnen - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="2" resultid="258" />
                    <RANKING place="3" resultid="259" />
                    <RANKING place="1" resultid="360" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="14" agemax="28" agemin="3" name="Offene Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="19" resultid="49" />
                    <RANKING place="51" resultid="50" />
                    <RANKING place="40" resultid="71" />
                    <RANKING place="21" resultid="142" />
                    <RANKING place="29" resultid="143" />
                    <RANKING place="41" resultid="144" />
                    <RANKING place="4" resultid="169" />
                    <RANKING place="3" resultid="258" />
                    <RANKING place="6" resultid="259" />
                    <RANKING place="13" resultid="260" />
                    <RANKING place="8" resultid="261" />
                    <RANKING place="14" resultid="263" />
                    <RANKING place="18" resultid="264" />
                    <RANKING place="27" resultid="266" />
                    <RANKING place="36" resultid="267" />
                    <RANKING place="60" resultid="268" />
                    <RANKING place="2" resultid="360" />
                    <RANKING place="10" resultid="361" />
                    <RANKING place="11" resultid="362" />
                    <RANKING place="22" resultid="363" />
                    <RANKING place="45" resultid="364" />
                    <RANKING place="43" resultid="365" />
                    <RANKING place="49" resultid="366" />
                    <RANKING place="58" resultid="367" />
                    <RANKING place="60" resultid="368" />
                    <RANKING place="26" resultid="518" />
                    <RANKING place="30" resultid="519" />
                    <RANKING place="34" resultid="520" />
                    <RANKING place="59" resultid="522" />
                    <RANKING place="63" resultid="524" />
                    <RANKING place="62" resultid="525" />
                    <RANKING place="24" resultid="692" />
                    <RANKING place="38" resultid="693" />
                    <RANKING place="5" resultid="748" />
                    <RANKING place="17" resultid="749" />
                    <RANKING place="19" resultid="750" />
                    <RANKING place="28" resultid="752" />
                    <RANKING place="37" resultid="753" />
                    <RANKING place="42" resultid="754" />
                    <RANKING place="50" resultid="755" />
                    <RANKING place="64" resultid="756" />
                    <RANKING place="7" resultid="915" />
                    <RANKING place="15" resultid="917" />
                    <RANKING place="12" resultid="918" />
                    <RANKING place="9" resultid="919" />
                    <RANKING place="16" resultid="921" />
                    <RANKING place="23" resultid="923" />
                    <RANKING place="35" resultid="924" />
                    <RANKING place="31" resultid="926" />
                    <RANKING place="44" resultid="927" />
                    <RANKING place="48" resultid="928" />
                    <RANKING place="57" resultid="929" />
                    <RANKING place="53" resultid="930" />
                    <RANKING place="47" resultid="931" />
                    <RANKING place="32" resultid="932" />
                    <RANKING place="1" resultid="1082" />
                    <RANKING place="25" resultid="1083" />
                    <RANKING place="33" resultid="1084" />
                    <RANKING place="39" resultid="1085" />
                    <RANKING place="46" resultid="1086" />
                    <RANKING place="52" resultid="1087" />
                    <RANKING place="54" resultid="1088" />
                    <RANKING place="56" resultid="1089" />
                    <RANKING place="55" resultid="1090" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="19" agemax="28" agemin="3" name="Offene internationale Wertung">
                  <RANKINGS>
                    <RANKING place="20" resultid="49" />
                    <RANKING place="57" resultid="50" />
                    <RANKING place="46" resultid="71" />
                    <RANKING place="22" resultid="142" />
                    <RANKING place="34" resultid="143" />
                    <RANKING place="47" resultid="144" />
                    <RANKING place="4" resultid="169" />
                    <RANKING place="3" resultid="258" />
                    <RANKING place="6" resultid="259" />
                    <RANKING place="14" resultid="260" />
                    <RANKING place="8" resultid="261" />
                    <RANKING place="15" resultid="263" />
                    <RANKING place="19" resultid="264" />
                    <RANKING place="32" resultid="266" />
                    <RANKING place="42" resultid="267" />
                    <RANKING place="66" resultid="268" />
                    <RANKING place="2" resultid="360" />
                    <RANKING place="10" resultid="361" />
                    <RANKING place="12" resultid="362" />
                    <RANKING place="23" resultid="363" />
                    <RANKING place="51" resultid="364" />
                    <RANKING place="49" resultid="365" />
                    <RANKING place="55" resultid="366" />
                    <RANKING place="64" resultid="367" />
                    <RANKING place="66" resultid="368" />
                    <RANKING place="11" resultid="408" />
                    <RANKING place="25" resultid="409" />
                    <RANKING place="27" resultid="410" />
                    <RANKING place="31" resultid="411" />
                    <RANKING place="30" resultid="518" />
                    <RANKING place="35" resultid="519" />
                    <RANKING place="39" resultid="520" />
                    <RANKING place="65" resultid="522" />
                    <RANKING place="69" resultid="524" />
                    <RANKING place="68" resultid="525" />
                    <RANKING place="29" resultid="665" />
                    <RANKING place="40" resultid="666" />
                    <RANKING place="26" resultid="692" />
                    <RANKING place="44" resultid="693" />
                    <RANKING place="5" resultid="748" />
                    <RANKING place="18" resultid="749" />
                    <RANKING place="20" resultid="750" />
                    <RANKING place="33" resultid="752" />
                    <RANKING place="43" resultid="753" />
                    <RANKING place="48" resultid="754" />
                    <RANKING place="56" resultid="755" />
                    <RANKING place="70" resultid="756" />
                    <RANKING place="7" resultid="915" />
                    <RANKING place="16" resultid="917" />
                    <RANKING place="13" resultid="918" />
                    <RANKING place="9" resultid="919" />
                    <RANKING place="17" resultid="921" />
                    <RANKING place="24" resultid="923" />
                    <RANKING place="41" resultid="924" />
                    <RANKING place="36" resultid="926" />
                    <RANKING place="50" resultid="927" />
                    <RANKING place="54" resultid="928" />
                    <RANKING place="63" resultid="929" />
                    <RANKING place="59" resultid="930" />
                    <RANKING place="53" resultid="931" />
                    <RANKING place="37" resultid="932" />
                    <RANKING place="1" resultid="1082" />
                    <RANKING place="28" resultid="1083" />
                    <RANKING place="38" resultid="1084" />
                    <RANKING place="45" resultid="1085" />
                    <RANKING place="52" resultid="1086" />
                    <RANKING place="58" resultid="1087" />
                    <RANKING place="60" resultid="1088" />
                    <RANKING place="62" resultid="1089" />
                    <RANKING place="61" resultid="1090" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15" agemax="44" agemin="29" name="Master A - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="4" resultid="170" />
                    <RANKING place="1" resultid="922" />
                    <RANKING place="3" resultid="925" />
                    <RANKING place="2" resultid="960" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="16" agemax="54" agemin="45" name="Master B - Süddeutsche Wertung" />
                <AGEGROUP agegroupid="17" agemax="-1" agemin="55" name="Master C - Süddeutsche Wertung" />
                <AGEGROUP agegroupid="18" agemax="-1" agemin="29" name="Offene internationale Wertung Master">
                  <RANKINGS>
                    <RANKING place="4" resultid="170" />
                    <RANKING place="1" resultid="922" />
                    <RANKING place="3" resultid="925" />
                    <RANKING place="2" resultid="960" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="17" number="17" gender="M" round="TIM">
              <SWIMSTYLE stroke="SURFACE" relaycount="1" distance="50" />
              <FEE value="500" currency="EUR" />
              <HEATS>
                <HEAT heatid="17001" number="1" />
                <HEAT heatid="17002" number="2" />
                <HEAT heatid="17003" number="3" />
                <HEAT heatid="17004" number="4" />
                <HEAT heatid="17005" number="5" />
                <HEAT heatid="17006" number="6" />
                <HEAT heatid="17007" number="7" />
                <HEAT heatid="17008" number="8" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="4" agemax="9" agemin="3" name="Jahrgang 2014 und jünger - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="2" resultid="57" />
                    <RANKING place="1" resultid="374" />
                    <RANKING place="3" resultid="535" />
                    <RANKING place="4" resultid="761" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="10" agemin="10" name="Jahrgang 2013 - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="2" resultid="56" />
                    <RANKING place="3" resultid="275" />
                    <RANKING place="1" resultid="276" />
                    <RANKING place="5" resultid="1093" />
                    <RANKING place="4" resultid="1094" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6" agemax="11" agemin="11" name="Jahrgang 2012 - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="2" resultid="55" />
                    <RANKING place="1" resultid="274" />
                    <RANKING place="3" resultid="373" />
                    <RANKING place="4" resultid="695" />
                    <RANKING place="5" resultid="943" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7" agemax="12" agemin="12" name="Jahrgang 2011 - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="2" resultid="273" />
                    <RANKING place="1" resultid="531" />
                    <RANKING place="3" resultid="759" />
                    <RANKING place="5" resultid="760" />
                    <RANKING place="4" resultid="1092" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8" agemax="13" agemin="13" name="Jahrgang 2010 - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="1" resultid="936" />
                    <RANKING place="2" resultid="938" />
                    <RANKING place="3" resultid="941" />
                    <RANKING place="4" resultid="942" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9" agemax="14" agemin="14" name="Jahrgang 2009 - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="1" resultid="53" />
                    <RANKING place="3" resultid="54" />
                    <RANKING place="2" resultid="372" />
                    <RANKING place="4" resultid="533" />
                    <RANKING place="5" resultid="940" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10" agemax="15" agemin="15" name="Jahrgang 2008 - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="3" resultid="52" />
                    <RANKING place="1" resultid="370" />
                    <RANKING place="2" resultid="935" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11" agemax="16" agemin="16" name="Jahrgang 2007 - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="1" resultid="758" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="12" agemax="17" agemin="17" name="Jahrgang 2006 - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="3" resultid="51" />
                    <RANKING place="2" resultid="527" />
                    <RANKING place="1" resultid="933" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="13" agemax="21" agemin="18" name="Junioren - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="2" resultid="269" />
                    <RANKING place="4" resultid="272" />
                    <RANKING place="1" resultid="526" />
                    <RANKING place="3" resultid="529" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="14" agemax="28" agemin="3" name="Offene Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="9" resultid="51" />
                    <RANKING place="13" resultid="52" />
                    <RANKING place="16" resultid="53" />
                    <RANKING place="20" resultid="54" />
                    <RANKING place="26" resultid="55" />
                    <RANKING place="30" resultid="56" />
                    <RANKING place="38" resultid="57" />
                    <RANKING place="4" resultid="269" />
                    <RANKING place="12" resultid="272" />
                    <RANKING place="19" resultid="273" />
                    <RANKING place="25" resultid="274" />
                    <RANKING place="31" resultid="275" />
                    <RANKING place="24" resultid="276" />
                    <RANKING place="6" resultid="369" />
                    <RANKING place="5" resultid="370" />
                    <RANKING place="17" resultid="372" />
                    <RANKING place="28" resultid="373" />
                    <RANKING place="33" resultid="374" />
                    <RANKING place="3" resultid="526" />
                    <RANKING place="7" resultid="527" />
                    <RANKING place="8" resultid="529" />
                    <RANKING place="15" resultid="531" />
                    <RANKING place="21" resultid="533" />
                    <RANKING place="40" resultid="535" />
                    <RANKING place="32" resultid="695" />
                    <RANKING place="2" resultid="757" />
                    <RANKING place="11" resultid="758" />
                    <RANKING place="27" resultid="759" />
                    <RANKING place="39" resultid="760" />
                    <RANKING place="41" resultid="761" />
                    <RANKING place="1" resultid="933" />
                    <RANKING place="10" resultid="935" />
                    <RANKING place="14" resultid="936" />
                    <RANKING place="18" resultid="938" />
                    <RANKING place="23" resultid="940" />
                    <RANKING place="22" resultid="941" />
                    <RANKING place="29" resultid="942" />
                    <RANKING place="37" resultid="943" />
                    <RANKING place="34" resultid="1092" />
                    <RANKING place="36" resultid="1093" />
                    <RANKING place="35" resultid="1094" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="19" agemax="28" agemin="3" name="Offene internationale Wertung">
                  <RANKINGS>
                    <RANKING place="12" resultid="51" />
                    <RANKING place="16" resultid="52" />
                    <RANKING place="20" resultid="53" />
                    <RANKING place="24" resultid="54" />
                    <RANKING place="30" resultid="55" />
                    <RANKING place="34" resultid="56" />
                    <RANKING place="42" resultid="57" />
                    <RANKING place="5" resultid="106" />
                    <RANKING place="11" resultid="107" />
                    <RANKING place="4" resultid="269" />
                    <RANKING place="15" resultid="272" />
                    <RANKING place="23" resultid="273" />
                    <RANKING place="29" resultid="274" />
                    <RANKING place="35" resultid="275" />
                    <RANKING place="28" resultid="276" />
                    <RANKING place="7" resultid="369" />
                    <RANKING place="6" resultid="370" />
                    <RANKING place="21" resultid="372" />
                    <RANKING place="32" resultid="373" />
                    <RANKING place="37" resultid="374" />
                    <RANKING place="9" resultid="412" />
                    <RANKING place="18" resultid="413" />
                    <RANKING place="3" resultid="526" />
                    <RANKING place="8" resultid="527" />
                    <RANKING place="10" resultid="529" />
                    <RANKING place="18" resultid="531" />
                    <RANKING place="25" resultid="533" />
                    <RANKING place="44" resultid="535" />
                    <RANKING place="36" resultid="695" />
                    <RANKING place="2" resultid="757" />
                    <RANKING place="14" resultid="758" />
                    <RANKING place="31" resultid="759" />
                    <RANKING place="43" resultid="760" />
                    <RANKING place="45" resultid="761" />
                    <RANKING place="1" resultid="933" />
                    <RANKING place="13" resultid="935" />
                    <RANKING place="17" resultid="936" />
                    <RANKING place="22" resultid="938" />
                    <RANKING place="27" resultid="940" />
                    <RANKING place="26" resultid="941" />
                    <RANKING place="33" resultid="942" />
                    <RANKING place="41" resultid="943" />
                    <RANKING place="38" resultid="1092" />
                    <RANKING place="40" resultid="1093" />
                    <RANKING place="39" resultid="1094" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15" agemax="44" agemin="29" name="Master A - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="1" resultid="171" />
                    <RANKING place="2" resultid="694" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="16" agemax="54" agemin="45" name="Master B - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="2" resultid="371" />
                    <RANKING place="1" resultid="934" />
                    <RANKING place="3" resultid="937" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="17" agemax="-1" agemin="55" name="Master C - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="1" resultid="121" />
                    <RANKING place="2" resultid="534" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="18" agemax="-1" agemin="29" name="Offene internationale Wertung Master">
                  <RANKINGS>
                    <RANKING place="4" resultid="121" />
                    <RANKING place="2" resultid="171" />
                    <RANKING place="5" resultid="371" />
                    <RANKING place="8" resultid="534" />
                    <RANKING place="7" resultid="694" />
                    <RANKING place="3" resultid="934" />
                    <RANKING place="6" resultid="937" />
                    <RANKING place="1" resultid="957" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="18" number="18" gender="F" round="TIM">
              <SWIMSTYLE stroke="BIFIN" relaycount="1" distance="50" />
              <FEE value="500" currency="EUR" />
              <HEATS>
                <HEAT heatid="18001" number="1" />
                <HEAT heatid="18002" number="2" />
                <HEAT heatid="18003" number="3" />
                <HEAT heatid="18004" number="4" />
                <HEAT heatid="18005" number="5" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="4" agemax="9" agemin="3" name="Jahrgang 2014 und jünger - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="2" resultid="251" />
                    <RANKING place="1" resultid="351" />
                    <RANKING place="4" resultid="499" />
                    <RANKING place="3" resultid="1063" />
                    <RANKING place="5" resultid="1064" />
                    <RANKING place="6" resultid="1065" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="10" agemin="10" name="Jahrgang 2013 - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="7" resultid="350" />
                    <RANKING place="4" resultid="898" />
                    <RANKING place="6" resultid="899" />
                    <RANKING place="1" resultid="1058" />
                    <RANKING place="2" resultid="1059" />
                    <RANKING place="5" resultid="1060" />
                    <RANKING place="8" resultid="1061" />
                    <RANKING place="3" resultid="1062" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6" agemax="11" agemin="11" name="Jahrgang 2012 - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="2" resultid="896" />
                    <RANKING place="1" resultid="897" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7" agemax="12" agemin="12" name="Jahrgang 2011 - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="3" resultid="349" />
                    <RANKING place="2" resultid="498" />
                    <RANKING place="1" resultid="1057" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8" agemax="13" agemin="13" name="Jahrgang 2010 - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="1" resultid="497" />
                    <RANKING place="2" resultid="1056" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9" agemax="14" agemin="14" name="Jahrgang 2009 - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="4" resultid="347" />
                    <RANKING place="1" resultid="890" />
                    <RANKING place="3" resultid="891" />
                    <RANKING place="2" resultid="892" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10" agemax="15" agemin="15" name="Jahrgang 2008 - Süddeutsche Wertung" />
                <AGEGROUP agegroupid="11" agemax="16" agemin="16" name="Jahrgang 2007 - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="1" resultid="140" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="12" agemax="17" agemin="17" name="Jahrgang 2006 - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="1" resultid="346" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="13" agemax="21" agemin="18" name="Juniorinnen - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="1" resultid="894" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="14" agemax="28" agemin="3" name="Offene Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="1" resultid="140" />
                    <RANKING place="24" resultid="251" />
                    <RANKING place="5" resultid="346" />
                    <RANKING place="8" resultid="347" />
                    <RANKING place="14" resultid="349" />
                    <RANKING place="21" resultid="350" />
                    <RANKING place="23" resultid="351" />
                    <RANKING place="7" resultid="497" />
                    <RANKING place="13" resultid="498" />
                    <RANKING place="26" resultid="499" />
                    <RANKING place="2" resultid="890" />
                    <RANKING place="4" resultid="891" />
                    <RANKING place="3" resultid="892" />
                    <RANKING place="6" resultid="894" />
                    <RANKING place="11" resultid="896" />
                    <RANKING place="10" resultid="897" />
                    <RANKING place="18" resultid="898" />
                    <RANKING place="20" resultid="899" />
                    <RANKING place="9" resultid="1056" />
                    <RANKING place="12" resultid="1057" />
                    <RANKING place="15" resultid="1058" />
                    <RANKING place="16" resultid="1059" />
                    <RANKING place="19" resultid="1060" />
                    <RANKING place="22" resultid="1061" />
                    <RANKING place="17" resultid="1062" />
                    <RANKING place="25" resultid="1063" />
                    <RANKING place="27" resultid="1064" />
                    <RANKING place="28" resultid="1065" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="19" agemax="28" agemin="3" name="Offene internationale Wertung">
                  <RANKINGS>
                    <RANKING place="1" resultid="103" />
                    <RANKING place="2" resultid="140" />
                    <RANKING place="25" resultid="251" />
                    <RANKING place="6" resultid="346" />
                    <RANKING place="9" resultid="347" />
                    <RANKING place="15" resultid="349" />
                    <RANKING place="22" resultid="350" />
                    <RANKING place="24" resultid="351" />
                    <RANKING place="8" resultid="497" />
                    <RANKING place="14" resultid="498" />
                    <RANKING place="27" resultid="499" />
                    <RANKING place="3" resultid="890" />
                    <RANKING place="5" resultid="891" />
                    <RANKING place="4" resultid="892" />
                    <RANKING place="7" resultid="894" />
                    <RANKING place="12" resultid="896" />
                    <RANKING place="11" resultid="897" />
                    <RANKING place="19" resultid="898" />
                    <RANKING place="21" resultid="899" />
                    <RANKING place="10" resultid="1056" />
                    <RANKING place="13" resultid="1057" />
                    <RANKING place="16" resultid="1058" />
                    <RANKING place="17" resultid="1059" />
                    <RANKING place="20" resultid="1060" />
                    <RANKING place="23" resultid="1061" />
                    <RANKING place="18" resultid="1062" />
                    <RANKING place="26" resultid="1063" />
                    <RANKING place="28" resultid="1064" />
                    <RANKING place="29" resultid="1065" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15" agemax="44" agemin="29" name="Master A - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="2" resultid="168" />
                    <RANKING place="1" resultid="893" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="16" agemax="54" agemin="45" name="Master B - Süddeutsche Wertung" />
                <AGEGROUP agegroupid="17" agemax="-1" agemin="55" name="Master C - Süddeutsche Wertung" />
                <AGEGROUP agegroupid="18" agemax="-1" agemin="29" name="Offene internationale Wertung Master">
                  <RANKINGS>
                    <RANKING place="2" resultid="168" />
                    <RANKING place="1" resultid="893" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="19" number="19" gender="M" round="TIM">
              <SWIMSTYLE stroke="BIFIN" relaycount="1" distance="50" />
              <FEE value="500" currency="EUR" />
              <HEATS>
                <HEAT heatid="19001" number="1" />
                <HEAT heatid="19002" number="2" />
                <HEAT heatid="19003" number="3" />
                <HEAT heatid="19004" number="4" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="4" agemax="9" agemin="3" name="Jahrgang 2014 und jünger - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="3" resultid="45" />
                    <RANKING place="1" resultid="355" />
                    <RANKING place="4" resultid="509" />
                    <RANKING place="2" resultid="904" />
                    <RANKING place="5" resultid="1069" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="10" agemin="10" name="Jahrgang 2013 - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="1" resultid="1067" />
                    <RANKING place="2" resultid="1068" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6" agemax="11" agemin="11" name="Jahrgang 2012 - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="1" resultid="354" />
                    <RANKING place="2" resultid="906" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7" agemax="12" agemin="12" name="Jahrgang 2011 - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="1" resultid="1066" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8" agemax="13" agemin="13" name="Jahrgang 2010 - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="3" resultid="506" />
                    <RANKING place="2" resultid="901" />
                    <RANKING place="1" resultid="902" />
                    <RANKING place="4" resultid="903" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9" agemax="14" agemin="14" name="Jahrgang 2009 - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="1" resultid="508" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10" agemax="15" agemin="15" name="Jahrgang 2008 - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="1" resultid="353" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11" agemax="16" agemin="16" name="Jahrgang 2007 - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="1" resultid="963" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="12" agemax="17" agemin="17" name="Jahrgang 2006 - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="2" resultid="252" />
                    <RANKING place="1" resultid="500" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="13" agemax="21" agemin="18" name="Junioren - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="3" resultid="501" />
                    <RANKING place="1" resultid="502" />
                    <RANKING place="2" resultid="504" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="14" agemax="28" agemin="3" name="Offene Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="19" resultid="45" />
                    <RANKING place="3" resultid="252" />
                    <RANKING place="1" resultid="352" />
                    <RANKING place="8" resultid="353" />
                    <RANKING place="13" resultid="354" />
                    <RANKING place="16" resultid="355" />
                    <RANKING place="2" resultid="500" />
                    <RANKING place="7" resultid="501" />
                    <RANKING place="4" resultid="502" />
                    <RANKING place="5" resultid="504" />
                    <RANKING place="11" resultid="506" />
                    <RANKING place="15" resultid="508" />
                    <RANKING place="22" resultid="509" />
                    <RANKING place="10" resultid="901" />
                    <RANKING place="9" resultid="902" />
                    <RANKING place="12" resultid="903" />
                    <RANKING place="17" resultid="904" />
                    <RANKING place="18" resultid="906" />
                    <RANKING place="6" resultid="963" />
                    <RANKING place="14" resultid="1066" />
                    <RANKING place="20" resultid="1067" />
                    <RANKING place="21" resultid="1068" />
                    <RANKING place="23" resultid="1069" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="19" agemax="28" agemin="3" name="Offene internationale Wertung">
                  <RANKINGS>
                    <RANKING place="19" resultid="45" />
                    <RANKING place="3" resultid="252" />
                    <RANKING place="1" resultid="352" />
                    <RANKING place="8" resultid="353" />
                    <RANKING place="13" resultid="354" />
                    <RANKING place="16" resultid="355" />
                    <RANKING place="2" resultid="500" />
                    <RANKING place="7" resultid="501" />
                    <RANKING place="4" resultid="502" />
                    <RANKING place="5" resultid="504" />
                    <RANKING place="11" resultid="506" />
                    <RANKING place="15" resultid="508" />
                    <RANKING place="22" resultid="509" />
                    <RANKING place="10" resultid="901" />
                    <RANKING place="9" resultid="902" />
                    <RANKING place="12" resultid="903" />
                    <RANKING place="17" resultid="904" />
                    <RANKING place="18" resultid="906" />
                    <RANKING place="6" resultid="963" />
                    <RANKING place="14" resultid="1066" />
                    <RANKING place="20" resultid="1067" />
                    <RANKING place="21" resultid="1068" />
                    <RANKING place="23" resultid="1069" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15" agemax="44" agemin="29" name="Master A - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="1" resultid="691" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="16" agemax="54" agemin="45" name="Master B - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="1" resultid="900" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="17" agemax="-1" agemin="55" name="Master C - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="1" resultid="120" />
                    <RANKING place="2" resultid="505" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="18" agemax="-1" agemin="29" name="Offene internationale Wertung Master">
                  <RANKINGS>
                    <RANKING place="2" resultid="120" />
                    <RANKING place="4" resultid="505" />
                    <RANKING place="5" resultid="691" />
                    <RANKING place="3" resultid="900" />
                    <RANKING place="1" resultid="956" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="20" number="20" gender="X" round="TIM">
              <SWIMSTYLE stroke="SURFACE" relaycount="1" distance="800" />
              <FEE value="500" currency="EUR" />
              <HEATS>
                <HEAT heatid="20001" number="1" />
                <HEAT heatid="20002" number="2" />
                <HEAT heatid="20003" number="3" />
                <HEAT heatid="20004" number="4" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="4" agemax="9" agemin="12" name="weiblich: Jahrgang 2014 und jünger - Süddeutsche Wertung" />
                <AGEGROUP agegroupid="5" agemax="10" agemin="12" name="weiblich: Jahrgang 2013 - Süddeutsche Wertung" />
                <AGEGROUP agegroupid="6" agemax="11" agemin="12" name="weiblich: Jahrgang 2012 - Süddeutsche Wertung" />
                <AGEGROUP agegroupid="7" agemax="12" agemin="12" name="weiblich: Jahrgang 2011 - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="1" resultid="379" />
                    <RANKING place="2" resultid="380" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8" agemax="13" agemin="13" name="weiblich: Jahrgang 2010 - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="2" resultid="538" />
                    <RANKING place="1" resultid="765" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9" agemax="14" agemin="14" name="weiblich: Jahrgang 2009 - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="1" resultid="949" />
                    <RANKING place="2" resultid="950" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10" agemax="15" agemin="15" name="weiblich: Jahrgang 2008 - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="1" resultid="767" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11" agemax="16" agemin="16" name="weiblich: Jahrgang 2007 - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="2" resultid="72" />
                    <RANKING place="1" resultid="145" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="12" agemax="17" agemin="17" name="weiblich: Jahrgang 2006 - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="1" resultid="696" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="13" agemax="21" agemin="18" name="Juniorinnen - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="1" resultid="1100" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="14" agemax="28" agemin="12" name="weiblich: Offene Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="9" resultid="60" />
                    <RANKING place="4" resultid="72" />
                    <RANKING place="2" resultid="145" />
                    <RANKING place="1" resultid="172" />
                    <RANKING place="10" resultid="379" />
                    <RANKING place="13" resultid="380" />
                    <RANKING place="12" resultid="538" />
                    <RANKING place="8" resultid="696" />
                    <RANKING place="11" resultid="765" />
                    <RANKING place="6" resultid="767" />
                    <RANKING place="3" resultid="949" />
                    <RANKING place="7" resultid="950" />
                    <RANKING place="5" resultid="1100" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="19" agemax="28" agemin="12" name="weiblich: Offene internationale Wertung">
                  <RANKINGS>
                    <RANKING place="10" resultid="60" />
                    <RANKING place="5" resultid="72" />
                    <RANKING place="2" resultid="109" />
                    <RANKING place="3" resultid="145" />
                    <RANKING place="1" resultid="172" />
                    <RANKING place="11" resultid="379" />
                    <RANKING place="14" resultid="380" />
                    <RANKING place="13" resultid="538" />
                    <RANKING place="9" resultid="696" />
                    <RANKING place="12" resultid="765" />
                    <RANKING place="7" resultid="767" />
                    <RANKING place="4" resultid="949" />
                    <RANKING place="8" resultid="950" />
                    <RANKING place="6" resultid="1100" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15" agemax="44" agemin="29" name="weiblich: Master A - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="1" resultid="961" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="16" agemax="54" agemin="45" name="weiblich: Master B - Süddeutsche Wertung" />
                <AGEGROUP agegroupid="17" agemax="-1" agemin="55" name="weiblich: Master C - Süddeutsche Wertung" />
                <AGEGROUP agegroupid="18" agemax="-1" agemin="29" name="weiblich: Offene internationale Wertung Master">
                  <RANKINGS>
                    <RANKING place="1" resultid="961" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="23" agemax="9" agemin="12" name="männlich: Jahrgang 2014 und jünger - Süddeutsche Wertung" />
                <AGEGROUP agegroupid="24" agemax="10" agemin="12" name="männlich: Jahrgang 2013 - Süddeutsche Wertung" />
                <AGEGROUP agegroupid="25" agemax="11" agemin="12" name="männlich: Jahrgang 2012 - Süddeutsche Wertung" />
                <AGEGROUP agegroupid="26" agemax="12" agemin="12" name="männlich: Jahrgang 2011 - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="1" resultid="378" />
                    <RANKING place="2" resultid="1099" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="27" agemax="13" agemin="13" name="männlich: Jahrgang 2010 - Süddeutsche Wertung" />
                <AGEGROUP agegroupid="28" agemax="14" agemin="14" name="männlich: Jahrgang 2009 - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="1" resultid="377" />
                    <RANKING place="2" resultid="951" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="29" agemax="15" agemin="15" name="männlich: Jahrgang 2008 - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="1" resultid="59" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="30" agemax="16" agemin="16" name="männlich: Jahrgang 2007 - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="1" resultid="766" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="31" agemax="17" agemin="17" name="männlich: Jahrgang 2006 - Süddeutsche Wertung" />
                <AGEGROUP agegroupid="32" agemax="21" agemin="18" name="Junioren - Süddeutsche Wertung" />
                <AGEGROUP agegroupid="33" agemax="28" agemin="12" name="männlich: Offene Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="1" resultid="59" />
                    <RANKING place="3" resultid="377" />
                    <RANKING place="5" resultid="378" />
                    <RANKING place="2" resultid="766" />
                    <RANKING place="4" resultid="951" />
                    <RANKING place="6" resultid="1099" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="38" agemax="28" agemin="12" name="männlich: Offene internationale Wertung">
                  <RANKINGS>
                    <RANKING place="2" resultid="59" />
                    <RANKING place="1" resultid="110" />
                    <RANKING place="4" resultid="377" />
                    <RANKING place="6" resultid="378" />
                    <RANKING place="3" resultid="766" />
                    <RANKING place="5" resultid="951" />
                    <RANKING place="7" resultid="1099" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="34" agemax="44" agemin="29" name="männlich: Master A - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="1" resultid="173" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="35" agemax="54" agemin="45" name="männlich: Master B - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="1" resultid="967" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="36" agemax="-1" agemin="55" name="männlich: Master C - Süddeutsche Wertung" />
                <AGEGROUP agegroupid="37" agemax="-1" agemin="29" name="männlich: Offene internationale Wertung Master">
                  <RANKINGS>
                    <RANKING place="1" resultid="173" />
                    <RANKING place="2" resultid="967" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="21" number="21" gender="F" round="TIM">
              <SWIMSTYLE stroke="IMMERSION" technique="DIVE" relaycount="1" distance="100" />
              <FEE value="500" currency="EUR" />
              <HEATS>
                <HEAT heatid="21001" number="1" />
                <HEAT heatid="21002" number="2" />
                <HEAT heatid="21003" number="3" />
                <HEAT heatid="21004" number="4" />
                <HEAT heatid="21005" number="5" />
                <HEAT heatid="21006" number="6" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="4" agemax="9" agemin="12" name="Jahrgang 2014 und jünger - Süddeutsche Wertung" />
                <AGEGROUP agegroupid="5" agemax="10" agemin="12" name="Jahrgang 2013 - Süddeutsche Wertung" />
                <AGEGROUP agegroupid="6" agemax="11" agemin="12" name="Jahrgang 2012 - Süddeutsche Wertung" />
                <AGEGROUP agegroupid="7" agemax="12" agemin="12" name="Jahrgang 2011 - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="1" resultid="129" />
                    <RANKING place="2" resultid="304" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8" agemax="13" agemin="13" name="Jahrgang 2010 - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="2" resultid="128" />
                    <RANKING place="4" resultid="714" />
                    <RANKING place="5" resultid="715" />
                    <RANKING place="1" resultid="810" />
                    <RANKING place="3" resultid="1017" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9" agemax="14" agemin="14" name="Jahrgang 2009 - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="2" resultid="195" />
                    <RANKING place="4" resultid="199" />
                    <RANKING place="3" resultid="303" />
                    <RANKING place="5" resultid="673" />
                    <RANKING place="1" resultid="809" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10" agemax="15" agemin="15" name="Jahrgang 2008 - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="1" resultid="198" />
                    <RANKING place="2" resultid="712" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11" agemax="16" agemin="16" name="Jahrgang 2007 - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="3" resultid="14" />
                    <RANKING place="2" resultid="64" />
                    <RANKING place="1" resultid="1016" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="12" agemax="17" agemin="17" name="Jahrgang 2006 - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="1" resultid="301" />
                    <RANKING place="4" resultid="672" />
                    <RANKING place="3" resultid="711" />
                    <RANKING place="2" resultid="808" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="13" agemax="21" agemin="18" name="Juniorinnen - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="1" resultid="127" />
                    <RANKING place="3" resultid="193" />
                    <RANKING place="4" resultid="194" />
                    <RANKING place="2" resultid="1014" />
                    <RANKING place="5" resultid="1015" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="14" agemax="28" agemin="12" name="Offene Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="29" resultid="14" />
                    <RANKING place="14" resultid="64" />
                    <RANKING place="1" resultid="127" />
                    <RANKING place="20" resultid="128" />
                    <RANKING place="26" resultid="129" />
                    <RANKING place="3" resultid="151" />
                    <RANKING place="5" resultid="193" />
                    <RANKING place="6" resultid="194" />
                    <RANKING place="15" resultid="195" />
                    <RANKING place="12" resultid="196" />
                    <RANKING place="17" resultid="198" />
                    <RANKING place="22" resultid="199" />
                    <RANKING place="9" resultid="301" />
                    <RANKING place="16" resultid="303" />
                    <RANKING place="28" resultid="304" />
                    <RANKING place="21" resultid="672" />
                    <RANKING place="27" resultid="673" />
                    <RANKING place="4" resultid="710" />
                    <RANKING place="18" resultid="711" />
                    <RANKING place="19" resultid="712" />
                    <RANKING place="24" resultid="714" />
                    <RANKING place="25" resultid="715" />
                    <RANKING place="11" resultid="808" />
                    <RANKING place="13" resultid="809" />
                    <RANKING place="10" resultid="810" />
                    <RANKING place="2" resultid="1014" />
                    <RANKING place="7" resultid="1015" />
                    <RANKING place="8" resultid="1016" />
                    <RANKING place="23" resultid="1017" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="19" agemax="28" agemin="12" name="Offene internationale Wertung">
                  <RANKINGS>
                    <RANKING place="33" resultid="14" />
                    <RANKING place="15" resultid="64" />
                    <RANKING place="9" resultid="81" />
                    <RANKING place="1" resultid="127" />
                    <RANKING place="23" resultid="128" />
                    <RANKING place="30" resultid="129" />
                    <RANKING place="3" resultid="151" />
                    <RANKING place="5" resultid="193" />
                    <RANKING place="6" resultid="194" />
                    <RANKING place="16" resultid="195" />
                    <RANKING place="13" resultid="196" />
                    <RANKING place="20" resultid="198" />
                    <RANKING place="26" resultid="199" />
                    <RANKING place="10" resultid="301" />
                    <RANKING place="18" resultid="303" />
                    <RANKING place="32" resultid="304" />
                    <RANKING place="17" resultid="387" />
                    <RANKING place="19" resultid="388" />
                    <RANKING place="25" resultid="389" />
                    <RANKING place="24" resultid="672" />
                    <RANKING place="31" resultid="673" />
                    <RANKING place="4" resultid="710" />
                    <RANKING place="21" resultid="711" />
                    <RANKING place="22" resultid="712" />
                    <RANKING place="28" resultid="714" />
                    <RANKING place="29" resultid="715" />
                    <RANKING place="12" resultid="808" />
                    <RANKING place="14" resultid="809" />
                    <RANKING place="11" resultid="810" />
                    <RANKING place="2" resultid="1014" />
                    <RANKING place="7" resultid="1015" />
                    <RANKING place="8" resultid="1016" />
                    <RANKING place="27" resultid="1017" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15" agemax="44" agemin="29" name="Master A - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="1" resultid="152" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="16" agemax="54" agemin="45" name="Master B - Süddeutsche Wertung" />
                <AGEGROUP agegroupid="17" agemax="-1" agemin="55" name="Master C - Süddeutsche Wertung" />
                <AGEGROUP agegroupid="18" agemax="-1" agemin="29" name="Offene internationale Wertung Master">
                  <RANKINGS>
                    <RANKING place="1" resultid="152" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="22" number="22" gender="M" round="TIM">
              <SWIMSTYLE stroke="IMMERSION" technique="DIVE" relaycount="1" distance="100" />
              <FEE value="500" currency="EUR" />
              <HEATS>
                <HEAT heatid="22001" number="1" />
                <HEAT heatid="22002" number="2" />
                <HEAT heatid="22003" number="3" />
                <HEAT heatid="22004" number="4" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="4" agemax="9" agemin="12" name="Jahrgang 2014 und jünger - Süddeutsche Wertung" />
                <AGEGROUP agegroupid="5" agemax="10" agemin="12" name="Jahrgang 2013 - Süddeutsche Wertung" />
                <AGEGROUP agegroupid="6" agemax="11" agemin="12" name="Jahrgang 2012 - Süddeutsche Wertung" />
                <AGEGROUP agegroupid="7" agemax="12" agemin="12" name="Jahrgang 2011 - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="1" resultid="203" />
                    <RANKING place="2" resultid="454" />
                    <RANKING place="3" resultid="718" />
                    <RANKING place="5" resultid="1018" />
                    <RANKING place="4" resultid="1019" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8" agemax="13" agemin="13" name="Jahrgang 2010 - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="2" resultid="453" />
                    <RANKING place="1" resultid="815" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9" agemax="14" agemin="14" name="Jahrgang 2009 - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="2" resultid="16" />
                    <RANKING place="1" resultid="305" />
                    <RANKING place="3" resultid="816" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10" agemax="15" agemin="15" name="Jahrgang 2008 - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="1" resultid="814" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11" agemax="16" agemin="16" name="Jahrgang 2007 - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="2" resultid="451" />
                    <RANKING place="1" resultid="717" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="12" agemax="17" agemin="17" name="Jahrgang 2006 - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="4" resultid="15" />
                    <RANKING place="2" resultid="201" />
                    <RANKING place="3" resultid="450" />
                    <RANKING place="1" resultid="811" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="13" agemax="21" agemin="18" name="Junioren - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="2" resultid="200" />
                    <RANKING place="1" resultid="446" />
                    <RANKING place="3" resultid="448" />
                    <RANKING place="4" resultid="449" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="14" agemax="28" agemin="12" name="Offene Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="11" resultid="15" />
                    <RANKING place="18" resultid="16" />
                    <RANKING place="4" resultid="200" />
                    <RANKING place="6" resultid="201" />
                    <RANKING place="15" resultid="203" />
                    <RANKING place="14" resultid="305" />
                    <RANKING place="2" resultid="446" />
                    <RANKING place="5" resultid="448" />
                    <RANKING place="7" resultid="449" />
                    <RANKING place="8" resultid="450" />
                    <RANKING place="10" resultid="451" />
                    <RANKING place="16" resultid="453" />
                    <RANKING place="17" resultid="454" />
                    <RANKING place="3" resultid="716" />
                    <RANKING place="9" resultid="717" />
                    <RANKING place="20" resultid="718" />
                    <RANKING place="1" resultid="811" />
                    <RANKING place="13" resultid="814" />
                    <RANKING place="12" resultid="815" />
                    <RANKING place="19" resultid="816" />
                    <RANKING place="22" resultid="1018" />
                    <RANKING place="21" resultid="1019" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="19" agemax="28" agemin="12" name="Offene internationale Wertung">
                  <RANKINGS>
                    <RANKING place="12" resultid="15" />
                    <RANKING place="20" resultid="16" />
                    <RANKING place="4" resultid="200" />
                    <RANKING place="7" resultid="201" />
                    <RANKING place="16" resultid="203" />
                    <RANKING place="15" resultid="305" />
                    <RANKING place="5" resultid="390" />
                    <RANKING place="18" resultid="391" />
                    <RANKING place="2" resultid="446" />
                    <RANKING place="6" resultid="448" />
                    <RANKING place="8" resultid="449" />
                    <RANKING place="9" resultid="450" />
                    <RANKING place="11" resultid="451" />
                    <RANKING place="17" resultid="453" />
                    <RANKING place="19" resultid="454" />
                    <RANKING place="3" resultid="716" />
                    <RANKING place="10" resultid="717" />
                    <RANKING place="22" resultid="718" />
                    <RANKING place="1" resultid="811" />
                    <RANKING place="14" resultid="814" />
                    <RANKING place="13" resultid="815" />
                    <RANKING place="21" resultid="816" />
                    <RANKING place="24" resultid="1018" />
                    <RANKING place="23" resultid="1019" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15" agemax="44" agemin="29" name="Master A - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="1" resultid="153" />
                    <RANKING place="2" resultid="674" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="16" agemax="54" agemin="45" name="Master B - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="1" resultid="812" />
                    <RANKING place="2" resultid="813" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="17" agemax="-1" agemin="55" name="Master C - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="1" resultid="452" />
                    <RANKING place="2" resultid="455" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="18" agemax="-1" agemin="29" name="Offene internationale Wertung Master">
                  <RANKINGS>
                    <RANKING place="1" resultid="153" />
                    <RANKING place="3" resultid="452" />
                    <RANKING place="6" resultid="455" />
                    <RANKING place="5" resultid="674" />
                    <RANKING place="2" resultid="812" />
                    <RANKING place="4" resultid="813" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="23" number="23" gender="F" round="TIM">
              <SWIMSTYLE stroke="FLY" technique="KICK" relaycount="1" distance="50" />
              <FEE value="500" currency="EUR" />
              <HEATS>
                <HEAT heatid="23001" number="1" />
                <HEAT heatid="23002" number="2" />
                <HEAT heatid="23003" number="3" />
                <HEAT heatid="23004" number="4" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="4" agemax="9" agemin="3" name="Jahrgang 2014 und jünger - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="1" resultid="357" />
                    <RANKING place="2" resultid="510" />
                    <RANKING place="4" resultid="746" />
                    <RANKING place="3" resultid="1072" />
                    <RANKING place="5" resultid="1078" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="10" agemin="10" name="Jahrgang 2013 - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="7" resultid="356" />
                    <RANKING place="5" resultid="907" />
                    <RANKING place="6" resultid="912" />
                    <RANKING place="1" resultid="1071" />
                    <RANKING place="4" resultid="1073" />
                    <RANKING place="2" resultid="1075" />
                    <RANKING place="3" resultid="1076" />
                    <RANKING place="8" resultid="1077" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6" agemax="11" agemin="11" name="Jahrgang 2012 - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="4" resultid="253" />
                    <RANKING place="2" resultid="254" />
                    <RANKING place="7" resultid="511" />
                    <RANKING place="9" resultid="514" />
                    <RANKING place="5" resultid="908" />
                    <RANKING place="3" resultid="909" />
                    <RANKING place="6" resultid="910" />
                    <RANKING place="8" resultid="911" />
                    <RANKING place="1" resultid="1070" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7" agemax="11" agemin="12" name="Jahrgang 2011 - Süddeutsche Wertung" />
                <AGEGROUP agegroupid="8" agemax="11" agemin="13" name="Jahrgang 2010 - Süddeutsche Wertung" />
                <AGEGROUP agegroupid="9" agemax="11" agemin="14" name="Jahrgang 2009 - Süddeutsche Wertung" />
                <AGEGROUP agegroupid="10" agemax="11" agemin="15" name="Jahrgang 2008 - Süddeutsche Wertung" />
                <AGEGROUP agegroupid="11" agemax="11" agemin="16" name="Jahrgang 2007 - Süddeutsche Wertung" />
                <AGEGROUP agegroupid="12" agemax="11" agemin="17" name="Jahrgang 2006 - Süddeutsche Wertung" />
                <AGEGROUP agegroupid="13" agemax="11" agemin="18" name="Juniorinnen - Süddeutsche Wertung" />
                <AGEGROUP agegroupid="14" agemax="11" agemin="3" name="Offene Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="4" resultid="253" />
                    <RANKING place="2" resultid="254" />
                    <RANKING place="20" resultid="356" />
                    <RANKING place="14" resultid="357" />
                    <RANKING place="15" resultid="510" />
                    <RANKING place="8" resultid="511" />
                    <RANKING place="17" resultid="514" />
                    <RANKING place="18" resultid="746" />
                    <RANKING place="13" resultid="907" />
                    <RANKING place="5" resultid="908" />
                    <RANKING place="3" resultid="909" />
                    <RANKING place="6" resultid="910" />
                    <RANKING place="10" resultid="911" />
                    <RANKING place="19" resultid="912" />
                    <RANKING place="1" resultid="1070" />
                    <RANKING place="7" resultid="1071" />
                    <RANKING place="16" resultid="1072" />
                    <RANKING place="12" resultid="1073" />
                    <RANKING place="9" resultid="1075" />
                    <RANKING place="11" resultid="1076" />
                    <RANKING place="22" resultid="1077" />
                    <RANKING place="21" resultid="1078" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="19" agemax="11" agemin="3" name="Offene internationale Wertung">
                  <RANKINGS>
                    <RANKING place="4" resultid="253" />
                    <RANKING place="2" resultid="254" />
                    <RANKING place="20" resultid="356" />
                    <RANKING place="14" resultid="357" />
                    <RANKING place="15" resultid="510" />
                    <RANKING place="8" resultid="511" />
                    <RANKING place="17" resultid="514" />
                    <RANKING place="18" resultid="746" />
                    <RANKING place="13" resultid="907" />
                    <RANKING place="5" resultid="908" />
                    <RANKING place="3" resultid="909" />
                    <RANKING place="6" resultid="910" />
                    <RANKING place="10" resultid="911" />
                    <RANKING place="19" resultid="912" />
                    <RANKING place="1" resultid="1070" />
                    <RANKING place="7" resultid="1071" />
                    <RANKING place="16" resultid="1072" />
                    <RANKING place="12" resultid="1073" />
                    <RANKING place="9" resultid="1075" />
                    <RANKING place="11" resultid="1076" />
                    <RANKING place="22" resultid="1077" />
                    <RANKING place="21" resultid="1078" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15" agemax="11" agemin="29" name="Master A - Süddeutsche Wertung" />
                <AGEGROUP agegroupid="16" agemax="11" agemin="45" name="Master B - Süddeutsche Wertung" />
                <AGEGROUP agegroupid="17" agemax="11" agemin="55" name="Master C - Süddeutsche Wertung" />
                <AGEGROUP agegroupid="18" agemax="11" agemin="29" name="Offene internationale Wertung Master" />
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="24" number="24" gender="M" round="TIM">
              <SWIMSTYLE stroke="FLY" technique="KICK" relaycount="1" distance="50" />
              <FEE value="500" currency="EUR" />
              <HEATS>
                <HEAT heatid="24001" number="1" />
                <HEAT heatid="24002" number="2" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="4" agemax="9" agemin="3" name="Jahrgang 2014 und jünger - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="2" resultid="48" />
                    <RANKING place="1" resultid="359" />
                    <RANKING place="4" resultid="515" />
                    <RANKING place="3" resultid="914" />
                    <RANKING place="5" resultid="1080" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="10" agemin="10" name="Jahrgang 2013 - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="2" resultid="47" />
                    <RANKING place="3" resultid="256" />
                    <RANKING place="1" resultid="257" />
                    <RANKING place="4" resultid="1081" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6" agemax="11" agemin="11" name="Jahrgang 2012 - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="3" resultid="46" />
                    <RANKING place="2" resultid="255" />
                    <RANKING place="1" resultid="358" />
                    <RANKING place="4" resultid="913" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7" agemax="11" agemin="12" name="Jahrgang 2011 - Süddeutsche Wertung" />
                <AGEGROUP agegroupid="8" agemax="11" agemin="13" name="Jahrgang 2010 - Süddeutsche Wertung" />
                <AGEGROUP agegroupid="9" agemax="11" agemin="14" name="Jahrgang 2009 - Süddeutsche Wertung" />
                <AGEGROUP agegroupid="10" agemax="11" agemin="15" name="Jahrgang 2008 - Süddeutsche Wertung" />
                <AGEGROUP agegroupid="11" agemax="11" agemin="16" name="Jahrgang 2007 - Süddeutsche Wertung" />
                <AGEGROUP agegroupid="12" agemax="11" agemin="17" name="Jahrgang 2006 - Süddeutsche Wertung" />
                <AGEGROUP agegroupid="13" agemax="11" agemin="18" name="Junioren - Süddeutsche Wertung" />
                <AGEGROUP agegroupid="14" agemax="11" agemin="3" name="Offene Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="3" resultid="46" />
                    <RANKING place="5" resultid="47" />
                    <RANKING place="9" resultid="48" />
                    <RANKING place="2" resultid="255" />
                    <RANKING place="7" resultid="256" />
                    <RANKING place="4" resultid="257" />
                    <RANKING place="1" resultid="358" />
                    <RANKING place="6" resultid="359" />
                    <RANKING place="11" resultid="515" />
                    <RANKING place="8" resultid="913" />
                    <RANKING place="10" resultid="914" />
                    <RANKING place="13" resultid="1080" />
                    <RANKING place="12" resultid="1081" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="19" agemax="11" agemin="3" name="Offene internationale Wertung">
                  <RANKINGS>
                    <RANKING place="3" resultid="46" />
                    <RANKING place="5" resultid="47" />
                    <RANKING place="9" resultid="48" />
                    <RANKING place="2" resultid="255" />
                    <RANKING place="7" resultid="256" />
                    <RANKING place="4" resultid="257" />
                    <RANKING place="1" resultid="358" />
                    <RANKING place="6" resultid="359" />
                    <RANKING place="11" resultid="515" />
                    <RANKING place="8" resultid="913" />
                    <RANKING place="10" resultid="914" />
                    <RANKING place="13" resultid="1080" />
                    <RANKING place="12" resultid="1081" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15" agemax="11" agemin="29" name="Master A - Süddeutsche Wertung" />
                <AGEGROUP agegroupid="16" agemax="11" agemin="45" name="Master B - Süddeutsche Wertung" />
                <AGEGROUP agegroupid="17" agemax="11" agemin="55" name="Master C - Süddeutsche Wertung" />
                <AGEGROUP agegroupid="18" agemax="11" agemin="29" name="Offene internationale Wertung Master" />
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="25" number="25" gender="F" round="TIM">
              <SWIMSTYLE stroke="SURFACE" relaycount="1" distance="400" />
              <FEE value="500" currency="EUR" />
              <HEATS>
                <HEAT heatid="25001" number="1" />
                <HEAT heatid="25002" number="2" />
                <HEAT heatid="25003" number="3" />
                <HEAT heatid="25004" number="4" />
                <HEAT heatid="25005" number="5" />
                <HEAT heatid="25006" number="6" />
                <HEAT heatid="25007" number="7" />
                <HEAT heatid="25008" number="8" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="4" agemax="9" agemin="10" name="Jahrgang 2014 und jünger - Süddeutsche Wertung" />
                <AGEGROUP agegroupid="5" agemax="10" agemin="10" name="Jahrgang 2013 - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="1" resultid="1035" />
                    <RANKING place="3" resultid="1039" />
                    <RANKING place="2" resultid="1040" />
                    <RANKING place="4" resultid="1041" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6" agemax="11" agemin="11" name="Jahrgang 2012 - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="2" resultid="222" />
                    <RANKING place="3" resultid="224" />
                    <RANKING place="5" resultid="735" />
                    <RANKING place="4" resultid="853" />
                    <RANKING place="6" resultid="854" />
                    <RANKING place="8" resultid="856" />
                    <RANKING place="7" resultid="858" />
                    <RANKING place="1" resultid="1036" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7" agemax="12" agemin="12" name="Jahrgang 2011 - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="4" resultid="223" />
                    <RANKING place="3" resultid="322" />
                    <RANKING place="7" resultid="323" />
                    <RANKING place="6" resultid="736" />
                    <RANKING place="1" resultid="852" />
                    <RANKING place="5" resultid="855" />
                    <RANKING place="2" resultid="1038" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8" agemax="13" agemin="13" name="Jahrgang 2010 - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="2" resultid="470" />
                    <RANKING place="3" resultid="733" />
                    <RANKING place="5" resultid="734" />
                    <RANKING place="1" resultid="847" />
                    <RANKING place="6" resultid="857" />
                    <RANKING place="4" resultid="1037" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9" agemax="14" agemin="14" name="Jahrgang 2009 - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="4" resultid="68" />
                    <RANKING place="1" resultid="218" />
                    <RANKING place="3" resultid="682" />
                    <RANKING place="2" resultid="849" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10" agemax="15" agemin="15" name="Jahrgang 2008 - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="1" resultid="731" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11" agemax="16" agemin="16" name="Jahrgang 2007 - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="3" resultid="31" />
                    <RANKING place="2" resultid="67" />
                    <RANKING place="1" resultid="136" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="12" agemax="17" agemin="17" name="Jahrgang 2006 - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="1" resultid="846" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="13" agemax="21" agemin="18" name="Juniorinnen - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="1" resultid="137" />
                    <RANKING place="4" resultid="216" />
                    <RANKING place="3" resultid="217" />
                    <RANKING place="2" resultid="321" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="14" agemax="28" agemin="10" name="Offene Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="8" resultid="30" />
                    <RANKING place="34" resultid="31" />
                    <RANKING place="9" resultid="67" />
                    <RANKING place="33" resultid="68" />
                    <RANKING place="7" resultid="136" />
                    <RANKING place="1" resultid="137" />
                    <RANKING place="2" resultid="158" />
                    <RANKING place="6" resultid="159" />
                    <RANKING place="5" resultid="216" />
                    <RANKING place="4" resultid="217" />
                    <RANKING place="10" resultid="218" />
                    <RANKING place="14" resultid="219" />
                    <RANKING place="18" resultid="222" />
                    <RANKING place="26" resultid="223" />
                    <RANKING place="24" resultid="224" />
                    <RANKING place="3" resultid="321" />
                    <RANKING place="22" resultid="322" />
                    <RANKING place="38" resultid="323" />
                    <RANKING place="17" resultid="470" />
                    <RANKING place="32" resultid="682" />
                    <RANKING place="13" resultid="731" />
                    <RANKING place="19" resultid="733" />
                    <RANKING place="30" resultid="734" />
                    <RANKING place="28" resultid="735" />
                    <RANKING place="35" resultid="736" />
                    <RANKING place="12" resultid="846" />
                    <RANKING place="11" resultid="847" />
                    <RANKING place="15" resultid="849" />
                    <RANKING place="20" resultid="852" />
                    <RANKING place="25" resultid="853" />
                    <RANKING place="29" resultid="854" />
                    <RANKING place="27" resultid="855" />
                    <RANKING place="39" resultid="856" />
                    <RANKING place="42" resultid="857" />
                    <RANKING place="31" resultid="858" />
                    <RANKING place="36" resultid="1035" />
                    <RANKING place="16" resultid="1036" />
                    <RANKING place="23" resultid="1037" />
                    <RANKING place="21" resultid="1038" />
                    <RANKING place="40" resultid="1039" />
                    <RANKING place="37" resultid="1040" />
                    <RANKING place="41" resultid="1041" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="19" agemax="28" agemin="10" name="Offene internationale Wertung">
                  <RANKINGS>
                    <RANKING place="10" resultid="30" />
                    <RANKING place="44" resultid="31" />
                    <RANKING place="11" resultid="67" />
                    <RANKING place="43" resultid="68" />
                    <RANKING place="1" resultid="89" />
                    <RANKING place="7" resultid="90" />
                    <RANKING place="23" resultid="92" />
                    <RANKING place="17" resultid="93" />
                    <RANKING place="9" resultid="136" />
                    <RANKING place="2" resultid="137" />
                    <RANKING place="3" resultid="158" />
                    <RANKING place="8" resultid="159" />
                    <RANKING place="6" resultid="216" />
                    <RANKING place="5" resultid="217" />
                    <RANKING place="12" resultid="218" />
                    <RANKING place="19" resultid="219" />
                    <RANKING place="27" resultid="222" />
                    <RANKING place="36" resultid="223" />
                    <RANKING place="34" resultid="224" />
                    <RANKING place="4" resultid="321" />
                    <RANKING place="32" resultid="322" />
                    <RANKING place="48" resultid="323" />
                    <RANKING place="16" resultid="397" />
                    <RANKING place="14" resultid="398" />
                    <RANKING place="25" resultid="399" />
                    <RANKING place="24" resultid="400" />
                    <RANKING place="26" resultid="470" />
                    <RANKING place="22" resultid="661" />
                    <RANKING place="30" resultid="662" />
                    <RANKING place="42" resultid="682" />
                    <RANKING place="18" resultid="731" />
                    <RANKING place="28" resultid="733" />
                    <RANKING place="40" resultid="734" />
                    <RANKING place="38" resultid="735" />
                    <RANKING place="45" resultid="736" />
                    <RANKING place="15" resultid="846" />
                    <RANKING place="13" resultid="847" />
                    <RANKING place="20" resultid="849" />
                    <RANKING place="29" resultid="852" />
                    <RANKING place="35" resultid="853" />
                    <RANKING place="39" resultid="854" />
                    <RANKING place="37" resultid="855" />
                    <RANKING place="49" resultid="856" />
                    <RANKING place="52" resultid="857" />
                    <RANKING place="41" resultid="858" />
                    <RANKING place="46" resultid="1035" />
                    <RANKING place="21" resultid="1036" />
                    <RANKING place="33" resultid="1037" />
                    <RANKING place="31" resultid="1038" />
                    <RANKING place="50" resultid="1039" />
                    <RANKING place="47" resultid="1040" />
                    <RANKING place="51" resultid="1041" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15" agemax="44" agemin="29" name="Master A - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="2" resultid="160" />
                    <RANKING place="1" resultid="848" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="16" agemax="54" agemin="45" name="Master B - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="1" resultid="469" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="17" agemax="-1" agemin="55" name="Master C - Süddeutsche Wertung" />
                <AGEGROUP agegroupid="18" agemax="-1" agemin="29" name="Offene internationale Wertung Master">
                  <RANKINGS>
                    <RANKING place="3" resultid="160" />
                    <RANKING place="1" resultid="469" />
                    <RANKING place="2" resultid="848" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="26" number="26" gender="M" round="TIM">
              <SWIMSTYLE stroke="SURFACE" relaycount="1" distance="400" />
              <FEE value="500" currency="EUR" />
              <HEATS>
                <HEAT heatid="26001" number="1" />
                <HEAT heatid="26002" number="2" />
                <HEAT heatid="26003" number="3" />
                <HEAT heatid="26004" number="4" />
                <HEAT heatid="26005" number="5" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="4" agemax="9" agemin="10" name="Jahrgang 2014 und jünger - Süddeutsche Wertung" />
                <AGEGROUP agegroupid="5" agemax="10" agemin="10" name="Jahrgang 2013 - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="2" resultid="36" />
                    <RANKING place="1" resultid="231" />
                    <RANKING place="5" resultid="232" />
                    <RANKING place="3" resultid="1042" />
                    <RANKING place="4" resultid="1043" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6" agemax="11" agemin="11" name="Jahrgang 2012 - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="4" resultid="37" />
                    <RANKING place="1" resultid="230" />
                    <RANKING place="2" resultid="328" />
                    <RANKING place="3" resultid="684" />
                    <RANKING place="5" resultid="859" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7" agemax="12" agemin="12" name="Jahrgang 2011 - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="1" resultid="229" />
                    <RANKING place="4" resultid="327" />
                    <RANKING place="6" resultid="738" />
                    <RANKING place="7" resultid="739" />
                    <RANKING place="2" resultid="976" />
                    <RANKING place="5" resultid="1044" />
                    <RANKING place="3" resultid="1045" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8" agemax="13" agemin="13" name="Jahrgang 2010 - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="1" resultid="861" />
                    <RANKING place="2" resultid="864" />
                    <RANKING place="3" resultid="865" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9" agemax="14" agemin="14" name="Jahrgang 2009 - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="2" resultid="34" />
                    <RANKING place="3" resultid="35" />
                    <RANKING place="1" resultid="325" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10" agemax="15" agemin="15" name="Jahrgang 2008 - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="1" resultid="324" />
                    <RANKING place="3" resultid="326" />
                    <RANKING place="2" resultid="862" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11" agemax="16" agemin="16" name="Jahrgang 2007 - Süddeutsche Wertung" />
                <AGEGROUP agegroupid="12" agemax="17" agemin="17" name="Jahrgang 2006 - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="3" resultid="33" />
                    <RANKING place="2" resultid="226" />
                    <RANKING place="1" resultid="860" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="13" agemax="21" agemin="18" name="Junioren - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="2" resultid="228" />
                    <RANKING place="1" resultid="471" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="14" agemax="28" agemin="10" name="Offene Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="6" resultid="33" />
                    <RANKING place="12" resultid="34" />
                    <RANKING place="15" resultid="35" />
                    <RANKING place="25" resultid="36" />
                    <RANKING place="28" resultid="37" />
                    <RANKING place="4" resultid="226" />
                    <RANKING place="5" resultid="228" />
                    <RANKING place="7" resultid="229" />
                    <RANKING place="16" resultid="230" />
                    <RANKING place="23" resultid="231" />
                    <RANKING place="29" resultid="232" />
                    <RANKING place="3" resultid="324" />
                    <RANKING place="9" resultid="325" />
                    <RANKING place="13" resultid="326" />
                    <RANKING place="20" resultid="327" />
                    <RANKING place="17" resultid="328" />
                    <RANKING place="2" resultid="471" />
                    <RANKING place="22" resultid="684" />
                    <RANKING place="24" resultid="738" />
                    <RANKING place="31" resultid="739" />
                    <RANKING place="30" resultid="859" />
                    <RANKING place="1" resultid="860" />
                    <RANKING place="8" resultid="861" />
                    <RANKING place="10" resultid="862" />
                    <RANKING place="14" resultid="864" />
                    <RANKING place="18" resultid="865" />
                    <RANKING place="11" resultid="976" />
                    <RANKING place="26" resultid="1042" />
                    <RANKING place="27" resultid="1043" />
                    <RANKING place="21" resultid="1044" />
                    <RANKING place="19" resultid="1045" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="19" agemax="28" agemin="10" name="Offene internationale Wertung">
                  <RANKINGS>
                    <RANKING place="7" resultid="33" />
                    <RANKING place="14" resultid="34" />
                    <RANKING place="17" resultid="35" />
                    <RANKING place="27" resultid="36" />
                    <RANKING place="30" resultid="37" />
                    <RANKING place="5" resultid="94" />
                    <RANKING place="4" resultid="226" />
                    <RANKING place="6" resultid="228" />
                    <RANKING place="9" resultid="229" />
                    <RANKING place="18" resultid="230" />
                    <RANKING place="25" resultid="231" />
                    <RANKING place="31" resultid="232" />
                    <RANKING place="3" resultid="324" />
                    <RANKING place="11" resultid="325" />
                    <RANKING place="15" resultid="326" />
                    <RANKING place="22" resultid="327" />
                    <RANKING place="19" resultid="328" />
                    <RANKING place="8" resultid="401" />
                    <RANKING place="2" resultid="471" />
                    <RANKING place="24" resultid="684" />
                    <RANKING place="26" resultid="738" />
                    <RANKING place="33" resultid="739" />
                    <RANKING place="32" resultid="859" />
                    <RANKING place="1" resultid="860" />
                    <RANKING place="10" resultid="861" />
                    <RANKING place="12" resultid="862" />
                    <RANKING place="16" resultid="864" />
                    <RANKING place="20" resultid="865" />
                    <RANKING place="13" resultid="976" />
                    <RANKING place="28" resultid="1042" />
                    <RANKING place="29" resultid="1043" />
                    <RANKING place="23" resultid="1044" />
                    <RANKING place="21" resultid="1045" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15" agemax="44" agemin="29" name="Master A - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="1" resultid="161" />
                    <RANKING place="2" resultid="683" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="16" agemax="54" agemin="45" name="Master B - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="1" resultid="968" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="17" agemax="-1" agemin="55" name="Master C - Süddeutsche Wertung" />
                <AGEGROUP agegroupid="18" agemax="-1" agemin="29" name="Offene internationale Wertung Master">
                  <RANKINGS>
                    <RANKING place="2" resultid="161" />
                    <RANKING place="4" resultid="683" />
                    <RANKING place="1" resultid="955" />
                    <RANKING place="3" resultid="968" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="27" number="27" gender="X" round="TIM">
              <SWIMSTYLE stroke="SURFACE" relaycount="4" distance="100" />
              <FEE value="800" currency="EUR" />
              <HEATS>
                <HEAT heatid="27001" number="1" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="2" agemax="11" agemin="3" name="Kategorie S3 - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="3" resultid="332" />
                    <RANKING place="1" resultid="870" />
                    <RANKING place="2" resultid="1049" />
                    <RANKING place="4" resultid="1103" />
                    <RANKING place="5" resultid="1104" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3" agemax="11" agemin="12" name="Kategorie S2 - Süddeutsche Wertung" />
                <AGEGROUP agegroupid="4" agemax="11" agemin="15" name="Kategorie S1 - Süddeutsche Wertung" />
                <AGEGROUP agegroupid="7" agemax="11" agemin="3" name="Offene Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="3" resultid="332" />
                    <RANKING place="1" resultid="870" />
                    <RANKING place="2" resultid="1049" />
                    <RANKING place="4" resultid="1103" />
                    <RANKING place="5" resultid="1104" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11" agemax="11" agemin="3" name="Offene internationale Wertung">
                  <RANKINGS>
                    <RANKING place="3" resultid="332" />
                    <RANKING place="1" resultid="870" />
                    <RANKING place="2" resultid="1049" />
                    <RANKING place="4" resultid="1103" />
                    <RANKING place="5" resultid="1104" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8" agemax="11" agemin="176" easy.ak="176" calculate="TOTAL" name="Masters A - Süddeutsche Wertung" />
                <AGEGROUP agegroupid="9" agemax="11" agemin="400" easy.ak="400" calculate="TOTAL" name="Masters B - Süddeutsche Wertung" />
                <AGEGROUP agegroupid="10" agemax="11" agemin="400" easy.ak="400" calculate="TOTAL" name="Offene internationale Wertung Master" />
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="28" number="28" gender="F" round="TIM">
              <SWIMSTYLE stroke="SURFACE" relaycount="4" distance="100" />
              <FEE value="800" currency="EUR" />
              <HEATS>
                <HEAT heatid="28001" number="1" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="2" agemax="11" agemin="12" name="Kategorie S3 - Süddeutsche Wertung" />
                <AGEGROUP agegroupid="3" agemax="14" agemin="12" name="Kategorie S2 - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="1" resultid="868" />
                    <RANKING place="2" resultid="869" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="17" agemin="15" name="Kategorie S1 - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="1" resultid="233" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7" agemax="123" agemin="12" name="Offene Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="3" resultid="233" />
                    <RANKING place="1" resultid="333" />
                    <RANKING place="2" resultid="868" />
                    <RANKING place="4" resultid="869" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11" agemax="123" agemin="12" name="Offene internationale Wertung">
                  <RANKINGS>
                    <RANKING place="1" resultid="96" />
                    <RANKING place="4" resultid="233" />
                    <RANKING place="2" resultid="333" />
                    <RANKING place="5" resultid="402" />
                    <RANKING place="3" resultid="868" />
                    <RANKING place="6" resultid="869" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8" agemax="-1" agemin="176" easy.ak="176" calculate="TOTAL" name="Masters A - Süddeutsche Wertung" />
                <AGEGROUP agegroupid="9" agemax="-1" agemin="400" easy.ak="400" calculate="TOTAL" name="Masters B - Süddeutsche Wertung" />
                <AGEGROUP agegroupid="10" agemax="-1" agemin="400" easy.ak="400" calculate="TOTAL" name="Offene internationale Wertung Master" />
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="29" number="29" gender="X" round="TIM">
              <SWIMSTYLE stroke="SURFACE" relaycount="4" distance="100" />
              <FEE value="800" currency="EUR" />
              <HEATS>
                <HEAT heatid="29001" number="1" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="2" agemax="11" agemin="12" name="Kategorie S3 - Süddeutsche Wertung" />
                <AGEGROUP agegroupid="3" agemax="14" agemin="12" name="Kategorie S2 - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="2" resultid="235" />
                    <RANKING place="1" resultid="872" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="17" agemin="15" name="Kategorie S1 - Süddeutsche Wertung" />
                <AGEGROUP agegroupid="7" agemax="123" agemin="12" name="Offene Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="3" resultid="235" />
                    <RANKING place="1" resultid="477" />
                    <RANKING place="2" resultid="872" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11" agemax="123" agemin="12" name="Offene internationale Wertung">
                  <RANKINGS>
                    <RANKING place="4" resultid="235" />
                    <RANKING place="1" resultid="477" />
                    <RANKING place="3" resultid="872" />
                    <RANKING place="2" resultid="975" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8" agemax="-1" agemin="176" easy.ak="176" calculate="TOTAL" name="Masters A - Süddeutsche Wertung" />
                <AGEGROUP agegroupid="9" agemax="-1" agemin="400" easy.ak="400" calculate="TOTAL" name="Masters B - Süddeutsche Wertung">
                  <RANKINGS>
                    <RANKING place="2" resultid="479" />
                    <RANKING place="1" resultid="871" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10" agemax="-1" agemin="400" easy.ak="400" calculate="TOTAL" name="Offene internationale Wertung Master">
                  <RANKINGS>
                    <RANKING place="2" resultid="479" />
                    <RANKING place="1" resultid="871" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
          </EVENTS>
        </SESSION>
      </SESSIONS>
      <CLUBS>
        <CLUB name="1. Chemnitzer Tauchverein e.V." nation="GER" region="20" code="0">
          <ATHLETES>
            <ATHLETE athleteid="90" birthdate="2008-01-01" gender="F" lastname="Franke" firstname="Jenny" license="0">
              <RESULTS>
                <RESULT resultid="381" eventid="1" swimtime="00:00:51.33" lane="4" heatid="1010" />
                <RESULT resultid="404" eventid="7" swimtime="00:00:21.65" lane="4" heatid="7003" />
                <RESULT resultid="392" eventid="11" swimtime="00:02:00.50" lane="5" heatid="11009">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:58.01" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="408" eventid="16" swimtime="00:00:23.28" lane="7" heatid="16010" />
                <RESULT resultid="387" eventid="21" swimtime="00:00:54.34" lane="6" heatid="21005" />
                <RESULT resultid="397" eventid="25" swimtime="00:04:21.51" lane="6" heatid="25007">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:00.10" />
                    <SPLIT distance="200" swimtime="00:02:08.40" />
                    <SPLIT distance="300" swimtime="00:03:17.03" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="91" birthdate="2007-01-01" gender="F" lastname="Ullrich" firstname="Johanna Hermine" license="0">
              <RESULTS>
                <RESULT resultid="382" eventid="1" swimtime="00:00:56.56" lane="1" heatid="1010" />
                <RESULT resultid="405" eventid="7" swimtime="00:00:24.39" lane="4" heatid="7002" />
                <RESULT resultid="393" eventid="11" swimtime="00:02:00.47" lane="3" heatid="11009">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:57.58" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="409" eventid="16" swimtime="00:00:25.88" lane="6" heatid="16009" />
                <RESULT resultid="388" eventid="21" swimtime="00:00:56.08" lane="2" heatid="21005" />
                <RESULT resultid="398" eventid="25" swimtime="00:04:18.47" lane="3" heatid="25006">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:59.23" />
                    <SPLIT distance="200" swimtime="00:02:06.32" />
                    <SPLIT distance="300" swimtime="00:03:14.47" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="92" birthdate="2010-01-01" gender="F" lastname="Schwarzer" firstname="Angelina Sophie" license="0">
              <RESULTS>
                <RESULT resultid="383" eventid="1" swimtime="00:00:58.14" lane="5" heatid="1008" />
                <RESULT resultid="414" eventid="9" swimtime="00:00:25.80" lane="6" heatid="9002" />
                <RESULT resultid="395" eventid="11" swimtime="00:02:12.98" lane="7" heatid="11007">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:03.39" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="410" eventid="16" swimtime="00:00:26.64" lane="2" heatid="16008" />
                <RESULT resultid="400" eventid="25" swimtime="00:04:54.49" lane="6" heatid="25005">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:06.49" />
                    <SPLIT distance="200" swimtime="00:02:24.17" />
                    <SPLIT distance="300" swimtime="00:03:43.33" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="93" birthdate="2011-01-01" gender="F" lastname="Nisch" firstname="Hanna Maria" license="0">
              <RESULTS>
                <RESULT resultid="384" eventid="1" swimtime="00:01:01.95" lane="4" heatid="1007" />
                <RESULT resultid="415" eventid="9" swimtime="00:00:27.03" lane="2" heatid="9002" />
                <RESULT resultid="394" eventid="11" swimtime="00:02:21.03" lane="8" heatid="11008">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:08.29" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="411" eventid="16" swimtime="00:00:27.35" lane="3" heatid="16007" />
                <RESULT resultid="389" eventid="21" swimtime="00:01:02.27" lane="2" heatid="21003" />
                <RESULT resultid="399" eventid="25" swimtime="00:05:06.46" lane="5" heatid="25005">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:13.38" />
                    <SPLIT distance="200" swimtime="00:02:34.49" />
                    <SPLIT distance="300" swimtime="00:03:54.15" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="94" birthdate="2006-01-01" gender="M" lastname="Lorenz" firstname="Emil" license="0">
              <RESULTS>
                <RESULT resultid="385" eventid="2" swimtime="00:00:43.18" lane="6" heatid="2008" />
                <RESULT resultid="406" eventid="8" swimtime="00:00:17.31" lane="6" heatid="8004" />
                <RESULT resultid="412" eventid="17" swimtime="00:00:20.07" lane="1" heatid="17008" />
                <RESULT resultid="390" eventid="22" swimtime="00:00:42.07" lane="1" heatid="22004" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="95" birthdate="2009-01-01" gender="M" lastname="Hans" firstname="Yannick" license="0">
              <RESULTS>
                <RESULT resultid="386" eventid="2" swimtime="00:00:54.77" lane="4" heatid="2005" />
                <RESULT resultid="407" eventid="8" swimtime="00:00:23.28" lane="2" heatid="8001" />
                <RESULT resultid="396" eventid="12" swimtime="00:02:00.54" lane="7" heatid="12006">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:58.44" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="413" eventid="17" swimtime="00:00:24.58" lane="8" heatid="17006" />
                <RESULT resultid="391" eventid="22" swimtime="00:00:59.47" lane="2" heatid="22002" />
                <RESULT resultid="401" eventid="26" swimtime="00:04:14.81" lane="5" heatid="26004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:56.94" />
                    <SPLIT distance="200" swimtime="00:02:04.58" />
                    <SPLIT distance="300" swimtime="00:03:12.37" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY number="1" gender="F" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="402" eventid="28" swimtime="00:03:49.53" lane="2" heatid="28001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:56.36" />
                    <SPLIT distance="200" swimtime="00:01:57.14" />
                    <SPLIT distance="300" swimtime="00:02:58.30" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="91" number="1" />
                    <RELAYPOSITION athleteid="92" number="2" />
                    <RELAYPOSITION athleteid="93" number="3" />
                    <RELAYPOSITION athleteid="90" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="2" gender="X" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="403" eventid="13" swimtime="00:01:35.04" lane="3" heatid="13001">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="95" number="1" />
                    <RELAYPOSITION athleteid="90" number="2" />
                    <RELAYPOSITION athleteid="92" number="3" />
                    <RELAYPOSITION athleteid="94" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB name="Aquanauten Karlsruhe-Durlach e.V." nation="GER" region="33" code="0">
          <ATHLETES>
            <ATHLETE athleteid="14" birthdate="2007-01-01" gender="F" lastname="Kirchner" firstname="Nia" license="0">
              <RESULTS>
                <RESULT resultid="62" eventid="1" swimtime="00:00:54.72" lane="7" heatid="1009" />
                <RESULT resultid="69" eventid="7" swimtime="00:00:23.10" lane="2" heatid="7002" />
                <RESULT resultid="65" eventid="15" swimtime="00:17:45.26" lane="8" heatid="15002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:04.16" />
                    <SPLIT distance="200" swimtime="00:02:14.39" />
                    <SPLIT distance="300" swimtime="00:03:26.49" />
                    <SPLIT distance="400" swimtime="00:04:38.45" />
                    <SPLIT distance="500" swimtime="00:05:50.65" />
                    <SPLIT distance="600" swimtime="00:07:05.03" />
                    <SPLIT distance="700" swimtime="00:08:17.45" />
                    <SPLIT distance="800" swimtime="00:09:29.96" />
                    <SPLIT distance="900" swimtime="00:10:44.57" />
                    <SPLIT distance="1000" swimtime="00:11:56.86" />
                    <SPLIT distance="1100" swimtime="00:13:10.44" />
                    <SPLIT distance="1200" swimtime="00:14:22.16" />
                    <SPLIT distance="1300" swimtime="00:15:34.67" />
                    <SPLIT distance="1400" swimtime="00:16:43.05" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="72" eventid="20" swimtime="00:08:43.54" lane="3" heatid="20003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:58.12" />
                    <SPLIT distance="200" swimtime="00:02:06.41" />
                    <SPLIT distance="300" swimtime="00:03:15.01" />
                    <SPLIT distance="400" swimtime="00:04:22.26" />
                    <SPLIT distance="500" swimtime="00:05:31.48" />
                    <SPLIT distance="600" swimtime="00:06:38.70" />
                    <SPLIT distance="700" swimtime="00:07:42.79" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="64" eventid="21" swimtime="00:00:52.96" lane="8" heatid="21005" />
                <RESULT resultid="67" eventid="25" swimtime="00:04:15.92" lane="7" heatid="25007">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:58.71" />
                    <SPLIT distance="200" swimtime="00:02:06.75" />
                    <SPLIT distance="300" swimtime="00:03:13.33" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="15" birthdate="2009-01-01" gender="F" lastname="Götte" firstname="Maja" license="0">
              <RESULTS>
                <RESULT resultid="63" eventid="1" swimtime="00:01:08.31" lane="3" heatid="1004" />
                <RESULT resultid="70" eventid="7" status="DSQ" swimtime="00:00:29.88" lane="3" heatid="7001" comment="falscher Start" />
                <RESULT resultid="66" eventid="11" swimtime="00:02:45.45" lane="8" heatid="11005">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:19.69" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="71" eventid="16" swimtime="00:00:30.53" lane="4" heatid="16004" />
                <RESULT resultid="68" eventid="25" swimtime="00:05:54.74" lane="7" heatid="25003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:19.33" />
                    <SPLIT distance="200" swimtime="00:02:53.02" />
                    <SPLIT distance="300" swimtime="00:04:28.03" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="Binger Tauchsportclub e.V." nation="GER" region="29" code="0">
          <ATHLETES>
            <ATHLETE athleteid="1" birthdate="2012-01-01" gender="M" lastname="Del Sordo" firstname="Ben" license="0">
              <RESULTS>
                <RESULT resultid="10" eventid="2" status="DSQ" swimtime="00:01:08.88" lane="2" heatid="2003" comment="falscher Start" />
                <RESULT resultid="1" eventid="4" swimtime="00:01:26.57" lane="6" heatid="4001" />
                <RESULT resultid="27" eventid="12" swimtime="00:02:40.95" lane="7" heatid="12003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:16.81" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="55" eventid="17" swimtime="00:00:31.01" lane="6" heatid="17003" />
                <RESULT resultid="46" eventid="24" swimtime="00:00:35.63" lane="4" heatid="24001" />
                <RESULT resultid="37" eventid="26" swimtime="00:06:27.47" lane="3" heatid="26001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:28.04" />
                    <SPLIT distance="200" swimtime="00:03:10.37" />
                    <SPLIT distance="300" swimtime="00:04:54.86" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="2" birthdate="2013-01-01" gender="M" lastname="Pieroth" firstname="Elias" license="0">
              <RESULTS>
                <RESULT resultid="11" eventid="2" swimtime="00:01:16.39" lane="1" heatid="2003" />
                <RESULT resultid="2" eventid="4" swimtime="00:01:24.42" lane="3" heatid="4001" />
                <RESULT resultid="26" eventid="12" swimtime="00:02:47.46" lane="5" heatid="12003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:20.93" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="56" eventid="17" swimtime="00:00:32.85" lane="1" heatid="17003" />
                <RESULT resultid="47" eventid="24" swimtime="00:00:36.33" lane="8" heatid="24002" />
                <RESULT resultid="36" eventid="26" swimtime="00:06:14.60" lane="5" heatid="26001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:31.74" />
                    <SPLIT distance="200" swimtime="00:03:09.28" />
                    <SPLIT distance="300" swimtime="00:04:47.95" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="3" birthdate="2014-01-01" gender="M" lastname="Gorsinsky" firstname="Felix" license="0">
              <RESULTS>
                <RESULT resultid="12" eventid="2" swimtime="00:01:30.51" lane="5" heatid="2001" />
                <RESULT resultid="3" eventid="4" swimtime="00:01:24.88" lane="2" heatid="4001" />
                <RESULT resultid="28" eventid="12" swimtime="00:03:06.06" lane="7" heatid="12002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:30.02" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="57" eventid="17" swimtime="00:00:40.60" lane="1" heatid="17002" />
                <RESULT resultid="45" eventid="19" swimtime="00:00:38.61" lane="4" heatid="19001" />
                <RESULT resultid="48" eventid="24" swimtime="00:00:42.17" lane="2" heatid="24001" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="4" birthdate="1997-01-01" gender="F" lastname="Walter" firstname="Lisa" license="0">
              <RESULTS>
                <RESULT resultid="4" eventid="1" swimtime="00:00:54.90" lane="3" heatid="1010" />
                <RESULT resultid="20" eventid="11" swimtime="00:02:00.29" lane="8" heatid="11010">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:57.91" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="19" eventid="15" swimtime="00:19:40.70" lane="5" heatid="15001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:11.00" />
                    <SPLIT distance="200" swimtime="00:02:29.06" />
                    <SPLIT distance="300" swimtime="00:03:48.21" />
                    <SPLIT distance="400" swimtime="00:05:07.65" />
                    <SPLIT distance="500" swimtime="00:06:28.05" />
                    <SPLIT distance="600" swimtime="00:07:46.86" />
                    <SPLIT distance="700" swimtime="00:09:07.27" />
                    <SPLIT distance="800" swimtime="00:10:27.02" />
                    <SPLIT distance="900" swimtime="00:11:47.31" />
                    <SPLIT distance="1000" swimtime="00:13:07.14" />
                    <SPLIT distance="1100" swimtime="00:14:28.69" />
                    <SPLIT distance="1200" swimtime="00:15:49.17" />
                    <SPLIT distance="1300" swimtime="00:17:08.33" />
                    <SPLIT distance="1400" swimtime="00:18:25.18" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="49" eventid="16" swimtime="00:00:25.55" lane="7" heatid="16009" />
                <RESULT resultid="60" eventid="20" swimtime="00:10:11.49" lane="2" heatid="20003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:10.24" />
                    <SPLIT distance="200" swimtime="00:02:27.06" />
                    <SPLIT distance="300" swimtime="00:03:44.71" />
                    <SPLIT distance="400" swimtime="00:05:03.16" />
                    <SPLIT distance="500" swimtime="00:06:21.09" />
                    <SPLIT distance="600" swimtime="00:07:39.11" />
                    <SPLIT distance="700" swimtime="00:08:56.34" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="30" eventid="25" swimtime="00:04:15.49" lane="5" heatid="25007">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:59.99" />
                    <SPLIT distance="200" swimtime="00:02:06.12" />
                    <SPLIT distance="300" swimtime="00:03:11.78" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="5" birthdate="2007-01-01" gender="F" lastname="Jöckel" firstname="Stella" license="0">
              <RESULTS>
                <RESULT resultid="5" eventid="1" swimtime="00:01:11.39" lane="7" heatid="1003" />
                <RESULT resultid="41" eventid="7" swimtime="00:00:33.64" lane="6" heatid="7001" />
                <RESULT resultid="21" eventid="11" status="DSQ" swimtime="00:02:48.97" lane="5" heatid="11004" comment="falsche Ausrüstung (Anzug) ">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:19.78" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="50" eventid="16" swimtime="00:00:33.67" lane="8" heatid="16004" />
                <RESULT resultid="14" eventid="21" swimtime="00:01:27.27" lane="5" heatid="21001" />
                <RESULT resultid="31" eventid="25" swimtime="00:05:57.01" lane="1" heatid="25002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:21.42" />
                    <SPLIT distance="200" swimtime="00:02:56.44" />
                    <SPLIT distance="300" swimtime="00:04:29.74" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="6" birthdate="2006-01-01" gender="M" lastname="Blaszczyk" firstname="Jan" license="0">
              <RESULTS>
                <RESULT resultid="6" eventid="2" swimtime="00:00:50.28" lane="5" heatid="2006" />
                <RESULT resultid="43" eventid="8" swimtime="00:00:20.01" lane="6" heatid="8001" />
                <RESULT resultid="23" eventid="12" swimtime="00:01:55.82" lane="6" heatid="12006">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:55.94" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="51" eventid="17" swimtime="00:00:21.94" lane="8" heatid="17007" />
                <RESULT resultid="15" eventid="22" swimtime="00:00:51.35" lane="5" heatid="22002" />
                <RESULT resultid="33" eventid="26" swimtime="00:04:13.42" lane="6" heatid="26004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:59.79" />
                    <SPLIT distance="200" swimtime="00:02:06.08" />
                    <SPLIT distance="300" swimtime="00:03:12.57" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="7" birthdate="2008-01-01" gender="M" lastname="Funke" firstname="Paul" license="0">
              <RESULTS>
                <RESULT resultid="7" eventid="2" swimtime="00:00:51.03" lane="3" heatid="2006" />
                <RESULT resultid="22" eventid="12" swimtime="00:01:56.31" lane="3" heatid="12006">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:56.18" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="17" eventid="15" swimtime="00:17:16.08" lane="2" heatid="15002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:04.46" />
                    <SPLIT distance="200" swimtime="00:02:14.89" />
                    <SPLIT distance="300" swimtime="00:03:25.11" />
                    <SPLIT distance="400" swimtime="00:04:35.12" />
                    <SPLIT distance="500" swimtime="00:05:44.68" />
                    <SPLIT distance="600" swimtime="00:06:54.48" />
                    <SPLIT distance="700" swimtime="00:08:03.69" />
                    <SPLIT distance="800" swimtime="00:09:14.11" />
                    <SPLIT distance="900" swimtime="00:10:23.29" />
                    <SPLIT distance="1000" swimtime="00:11:32.77" />
                    <SPLIT distance="1100" swimtime="00:12:42.25" />
                    <SPLIT distance="1200" swimtime="00:13:52.27" />
                    <SPLIT distance="1300" swimtime="00:15:01.70" />
                    <SPLIT distance="1400" swimtime="00:16:09.84" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="52" eventid="17" swimtime="00:00:23.30" lane="3" heatid="17006" />
                <RESULT resultid="59" eventid="20" swimtime="00:08:45.38" lane="8" heatid="20004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:01.05" />
                    <SPLIT distance="200" swimtime="00:02:06.17" />
                    <SPLIT distance="300" swimtime="00:03:13.16" />
                    <SPLIT distance="400" swimtime="00:04:21.16" />
                    <SPLIT distance="500" swimtime="00:05:29.35" />
                    <SPLIT distance="600" swimtime="00:06:37.23" />
                    <SPLIT distance="700" swimtime="00:07:42.68" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="32" eventid="26" status="DNS" swimtime="00:00:00.00" lane="1" heatid="26005" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="8" birthdate="2009-01-01" gender="M" lastname="Moritz" firstname="Silas" license="0">
              <RESULTS>
                <RESULT resultid="8" eventid="2" swimtime="00:00:54.67" lane="5" heatid="2005" />
                <RESULT resultid="42" eventid="8" swimtime="00:00:22.51" lane="1" heatid="8002" />
                <RESULT resultid="24" eventid="12" swimtime="00:02:07.98" lane="8" heatid="12006">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:02.02" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="18" eventid="15" status="DNS" swimtime="00:00:00.00" lane="1" heatid="15002" />
                <RESULT resultid="53" eventid="17" swimtime="00:00:25.18" lane="1" heatid="17006" />
                <RESULT resultid="61" eventid="20" status="DNS" swimtime="00:00:00.00" lane="1" heatid="20003" />
                <RESULT resultid="34" eventid="26" swimtime="00:04:38.19" lane="1" heatid="26004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:05.49" />
                    <SPLIT distance="200" swimtime="00:02:18.08" />
                    <SPLIT distance="300" swimtime="00:03:33.09" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="9" birthdate="2009-01-01" gender="M" lastname="Blaszczyk" firstname="Leonard" license="0">
              <RESULTS>
                <RESULT resultid="9" eventid="2" swimtime="00:00:59.45" lane="5" heatid="2004" />
                <RESULT resultid="44" eventid="8" swimtime="00:00:25.32" lane="7" heatid="8001" />
                <RESULT resultid="25" eventid="12" swimtime="00:02:12.61" lane="8" heatid="12005">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:01.44" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="54" eventid="17" swimtime="00:00:27.35" lane="8" heatid="17005" />
                <RESULT resultid="16" eventid="22" swimtime="00:01:06.10" lane="8" heatid="22002" />
                <RESULT resultid="35" eventid="26" swimtime="00:05:08.09" lane="5" heatid="26003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:07.69" />
                    <SPLIT distance="200" swimtime="00:02:28.19" />
                    <SPLIT distance="300" swimtime="00:03:51.62" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="10" birthdate="2017-01-01" gender="M" lastname="Pieroth" firstname="Milan" license="0">
              <RESULTS>
                <RESULT resultid="13" eventid="2" status="DSQ" swimtime="00:00:00.00" lane="3" heatid="2001" comment="Aufgegeben nach 20 m" />
                <RESULT resultid="29" eventid="12" status="DNS" swimtime="00:00:00.00" lane="5" heatid="12001" />
                <RESULT resultid="58" eventid="17" status="DNS" swimtime="00:00:00.00" lane="3" heatid="17001" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY number="1" gender="M" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="38" eventid="27" status="DNS" swimtime="00:00:00.00" lane="2" heatid="27001">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1" number="1" />
                    <RELAYPOSITION athleteid="2" number="2" />
                    <RELAYPOSITION athleteid="3" number="3" />
                    <RELAYPOSITION athleteid="10" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" gender="M" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="39" eventid="29" status="DNS" swimtime="00:00:00.00" lane="3" heatid="29001">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="6" number="1" />
                    <RELAYPOSITION athleteid="9" number="2" />
                    <RELAYPOSITION athleteid="8" number="3" />
                    <RELAYPOSITION athleteid="7" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" gender="X" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="40" eventid="13" swimtime="00:01:46.43" lane="6" heatid="13001">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4" number="1" />
                    <RELAYPOSITION athleteid="5" number="2" />
                    <RELAYPOSITION athleteid="6" number="3" />
                    <RELAYPOSITION athleteid="9" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB name="SC DHfK Leipzig Flossenschwimmen" nation="GER" region="20" code="0">
          <ATHLETES>
            <ATHLETE athleteid="16" birthdate="2008-01-01" gender="F" lastname="Kulchytska" firstname="Polina" license="0">
              <RESULTS>
                <RESULT resultid="73" eventid="1" swimtime="00:00:49.80" lane="4" heatid="1011" />
                <RESULT resultid="109" eventid="20" swimtime="00:08:08.66" lane="5" heatid="20004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:57.52" />
                    <SPLIT distance="200" swimtime="00:01:59.78" />
                    <SPLIT distance="300" swimtime="00:03:02.42" />
                    <SPLIT distance="400" swimtime="00:04:04.97" />
                    <SPLIT distance="500" swimtime="00:05:06.35" />
                    <SPLIT distance="600" swimtime="00:06:07.97" />
                    <SPLIT distance="700" swimtime="00:07:09.18" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="81" eventid="21" swimtime="00:00:46.91" lane="8" heatid="21006" />
                <RESULT resultid="90" eventid="25" swimtime="00:03:58.46" lane="3" heatid="25008">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:56.67" />
                    <SPLIT distance="200" swimtime="00:01:59.55" />
                    <SPLIT distance="300" swimtime="00:03:00.18" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="18" birthdate="2008-01-01" gender="F" lastname="Säbisch" firstname="Kyra" license="0">
              <RESULTS>
                <RESULT resultid="75" eventid="1" swimtime="00:00:52.15" lane="4" heatid="1009" />
                <RESULT resultid="99" eventid="7" swimtime="00:00:21.08" lane="2" heatid="7004" />
                <RESULT resultid="83" eventid="11" swimtime="00:02:00.13" lane="6" heatid="11008">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:55.88" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="104" eventid="16" status="DSQ" swimtime="00:00:23.33" lane="4" heatid="16010" comment="15m nach Start übertaucht" />
                <RESULT resultid="93" eventid="25" swimtime="00:04:26.72" lane="2" heatid="25005">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:58.42" />
                    <SPLIT distance="200" swimtime="00:02:06.51" />
                    <SPLIT distance="300" swimtime="00:03:17.59" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="19" birthdate="2010-01-01" gender="F" lastname="Horenok" firstname="Polina" license="0">
              <RESULTS>
                <RESULT resultid="76" eventid="1" swimtime="00:00:59.58" lane="7" heatid="1008" />
                <RESULT resultid="84" eventid="11" swimtime="00:02:15.30" lane="1" heatid="11007">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:05.90" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="105" eventid="16" status="DSQ" swimtime="00:00:26.09" lane="7" heatid="16008" comment="Tauchzüge (bei 45-50m)" />
                <RESULT resultid="92" eventid="25" swimtime="00:04:53.20" lane="1" heatid="25006">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:07.68" />
                    <SPLIT distance="200" swimtime="00:02:25.84" />
                    <SPLIT distance="300" swimtime="00:03:43.21" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="20" birthdate="2001-01-01" gender="M" lastname="Mörstedt" firstname="Justus" license="0">
              <RESULTS>
                <RESULT resultid="77" eventid="2" swimtime="00:00:35.00" lane="4" heatid="2008" />
                <RESULT resultid="95" eventid="6" swimtime="00:02:52.21" lane="4" heatid="6002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:39.93" />
                    <SPLIT distance="200" swimtime="00:01:22.69" />
                    <SPLIT distance="300" swimtime="00:02:07.00" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="85" eventid="12" swimtime="00:01:23.56" lane="4" heatid="12007">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:40.90" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="21" birthdate="2007-01-01" gender="M" lastname="Schoodt" firstname="Ben Joseph" license="0">
              <RESULTS>
                <RESULT resultid="78" eventid="2" swimtime="00:00:43.42" lane="5" heatid="2007" />
                <RESULT resultid="101" eventid="8" swimtime="00:00:17.84" lane="1" heatid="8004" />
                <RESULT resultid="86" eventid="12" swimtime="00:01:42.52" lane="3" heatid="12007">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:49.35" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="106" eventid="17" swimtime="00:00:19.30" lane="3" heatid="17008" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="22" birthdate="2008-01-01" gender="M" lastname="Berger" firstname="Alex Michael" license="0">
              <RESULTS>
                <RESULT resultid="79" eventid="2" swimtime="00:00:47.31" lane="7" heatid="2007" />
                <RESULT resultid="87" eventid="12" swimtime="00:01:47.80" lane="8" heatid="12007">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:51.28" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="107" eventid="17" swimtime="00:00:21.19" lane="7" heatid="17007" />
                <RESULT resultid="110" eventid="20" swimtime="00:08:25.48" lane="2" heatid="20004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:57.98" />
                    <SPLIT distance="200" swimtime="00:02:02.47" />
                    <SPLIT distance="300" swimtime="00:03:07.48" />
                    <SPLIT distance="400" swimtime="00:04:13.82" />
                    <SPLIT distance="500" swimtime="00:05:18.82" />
                    <SPLIT distance="600" swimtime="00:06:23.99" />
                    <SPLIT distance="700" swimtime="00:07:27.77" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="23" birthdate="2009-01-01" gender="M" lastname="Batiuk" firstname="Mykyta" license="0">
              <RESULTS>
                <RESULT resultid="80" eventid="2" swimtime="00:00:45.12" lane="4" heatid="2006" />
                <RESULT resultid="102" eventid="8" swimtime="00:00:17.91" lane="4" heatid="8002" />
                <RESULT resultid="88" eventid="12" swimtime="00:01:46.52" lane="6" heatid="12005">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:50.05" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="108" eventid="17" status="DSQ" swimtime="00:00:20.39" lane="1" heatid="17007" comment="15m nach Start übertaucht" />
                <RESULT resultid="94" eventid="26" swimtime="00:04:05.16" lane="8" heatid="26005">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:54.55" />
                    <SPLIT distance="200" swimtime="00:02:00.01" />
                    <SPLIT distance="300" swimtime="00:03:05.35" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="24" birthdate="2008-01-01" gender="F" lastname="Horenok" firstname="Maiia" license="0">
              <RESULTS>
                <RESULT resultid="103" eventid="18" swimtime="00:00:24.92" lane="5" heatid="18005" />
                <RESULT resultid="89" eventid="25" swimtime="00:03:41.24" lane="5" heatid="25008">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:52.08" />
                    <SPLIT distance="200" swimtime="00:01:48.28" />
                    <SPLIT distance="300" swimtime="00:02:46.23" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="28" birthdate="1977-01-01" gender="M" lastname="Nehrdich" firstname="Thomas" license="0">
              <RESULTS>
                <RESULT resultid="953" eventid="2" swimtime="00:00:46.22" lane="8" heatid="2007" />
                <RESULT resultid="952" eventid="4" swimtime="00:00:53.94" lane="3" heatid="4003" />
                <RESULT resultid="954" eventid="12" swimtime="00:01:49.62" lane="4" heatid="12006">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:54.03" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="957" eventid="17" swimtime="00:00:20.48" lane="4" heatid="17007" />
                <RESULT resultid="956" eventid="19" swimtime="00:00:24.14" lane="3" heatid="19004" />
                <RESULT resultid="955" eventid="26" swimtime="00:03:54.39" lane="7" heatid="26005">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:52.56" />
                    <SPLIT distance="200" swimtime="00:01:53.36" />
                    <SPLIT distance="300" swimtime="00:02:56.93" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY number="1" gender="F" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="96" eventid="28" swimtime="00:03:26.90" lane="5" heatid="28001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:50.81" />
                    <SPLIT distance="200" swimtime="00:01:49.78" />
                    <SPLIT distance="300" swimtime="00:02:42.06" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="16" number="1" />
                    <RELAYPOSITION athleteid="19" number="2" />
                    <RELAYPOSITION athleteid="18" number="3" />
                    <RELAYPOSITION athleteid="24" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" gender="X" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="98" eventid="13" swimtime="00:01:25.38" lane="5" heatid="13003">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="21" number="1" />
                    <RELAYPOSITION athleteid="23" number="2" />
                    <RELAYPOSITION athleteid="18" number="3" />
                    <RELAYPOSITION athleteid="16" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" gender="M" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="975" eventid="29" swimtime="00:03:05.34" lane="4" heatid="29001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:46.59" />
                    <SPLIT distance="200" swimtime="00:01:34.04" />
                    <SPLIT distance="300" swimtime="00:02:23.29" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="28" number="1" />
                    <RELAYPOSITION athleteid="23" number="2" />
                    <RELAYPOSITION athleteid="22" number="3" />
                    <RELAYPOSITION athleteid="21" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB name="SC Riesa e.V. Sekt. FS" nation="GER" region="20" code="0">
          <ATHLETES>
            <ATHLETE athleteid="159" birthdate="2010-01-01" gender="F" lastname="Berger" firstname="Lene" license="0">
              <RESULTS>
                <RESULT resultid="657" eventid="1" status="DSQ" swimtime="00:00:59.29" lane="4" heatid="1005" comment="falscher Start" />
                <RESULT resultid="659" eventid="11" swimtime="00:02:21.44" lane="8" heatid="11007">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:03.98" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="665" eventid="16" swimtime="00:00:27.17" lane="5" heatid="16005" />
                <RESULT resultid="661" eventid="25" swimtime="00:04:51.98" lane="8" heatid="25003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:06.15" />
                    <SPLIT distance="200" swimtime="00:02:21.43" />
                    <SPLIT distance="300" swimtime="00:03:39.24" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="160" birthdate="2011-01-01" gender="F" lastname="Hönisch" firstname="Ida" license="0">
              <RESULTS>
                <RESULT resultid="658" eventid="1" swimtime="00:01:03.68" lane="6" heatid="1005" />
                <RESULT resultid="660" eventid="11" swimtime="00:02:27.84" lane="7" heatid="11005">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:08.26" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="666" eventid="16" swimtime="00:00:29.12" lane="2" heatid="16005" />
                <RESULT resultid="662" eventid="25" swimtime="00:05:14.53" lane="3" heatid="25002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:06.47" />
                    <SPLIT distance="200" swimtime="00:02:24.71" />
                    <SPLIT distance="300" swimtime="00:03:45.24" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="161" birthdate="2006-01-01" gender="M" lastname="Loßner" firstname="Niklas" license="0">
              <RESULTS>
                <RESULT resultid="663" eventid="6" swimtime="00:03:18.85" lane="3" heatid="6002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:44.44" />
                    <SPLIT distance="200" swimtime="00:01:34.47" />
                    <SPLIT distance="300" swimtime="00:02:27.35" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="664" eventid="8" swimtime="00:00:15.10" lane="4" heatid="8004" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="SG Finswimming Jena" nation="GER" region="35" code="0">
          <ATHLETES>
            <ATHLETE athleteid="162" birthdate="2006-01-01" gender="F" lastname="Fabian" firstname="Lareen" license="0">
              <RESULTS>
                <RESULT resultid="667" eventid="1" swimtime="00:00:56.85" lane="3" heatid="1009" />
                <RESULT resultid="688" eventid="7" swimtime="00:00:23.55" lane="1" heatid="7003" />
                <RESULT resultid="677" eventid="11" swimtime="00:02:10.35" lane="3" heatid="11008">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:02.23" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="692" eventid="16" swimtime="00:00:26.01" lane="5" heatid="16008" />
                <RESULT resultid="696" eventid="20" swimtime="00:10:10.06" lane="4" heatid="20002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:03.43" />
                    <SPLIT distance="200" swimtime="00:02:18.44" />
                    <SPLIT distance="300" swimtime="00:03:36.11" />
                    <SPLIT distance="400" swimtime="00:04:55.25" />
                    <SPLIT distance="500" swimtime="00:06:15.32" />
                    <SPLIT distance="600" swimtime="00:07:35.16" />
                    <SPLIT distance="700" swimtime="00:08:54.77" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="672" eventid="21" swimtime="00:01:00.48" lane="3" heatid="21003" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="163" birthdate="2009-01-01" gender="F" lastname="Steininger" firstname="Magda" license="0">
              <RESULTS>
                <RESULT resultid="668" eventid="1" swimtime="00:00:57.22" lane="1" heatid="1008" />
                <RESULT resultid="689" eventid="7" swimtime="00:00:24.53" lane="7" heatid="7002" />
                <RESULT resultid="676" eventid="11" swimtime="00:02:15.21" lane="1" heatid="11009">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:02.97" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="164" birthdate="2009-01-01" gender="F" lastname="Fabian" firstname="Ileen" license="0">
              <RESULTS>
                <RESULT resultid="669" eventid="1" swimtime="00:01:10.22" lane="8" heatid="1005" />
                <RESULT resultid="678" eventid="11" status="DSQ" swimtime="00:02:41.22" lane="1" heatid="11005" comment="falscher Start">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:11.92" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="693" eventid="16" swimtime="00:00:30.03" lane="3" heatid="16005" />
                <RESULT resultid="673" eventid="21" swimtime="00:01:18.25" lane="4" heatid="21001" />
                <RESULT resultid="682" eventid="25" swimtime="00:05:48.09" lane="3" heatid="25005">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:15.03" />
                    <SPLIT distance="200" swimtime="00:02:44.76" />
                    <SPLIT distance="300" swimtime="00:04:17.60" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="166" birthdate="2012-01-01" gender="M" lastname="Gerbach" firstname="Linus" license="0">
              <RESULTS>
                <RESULT resultid="671" eventid="2" swimtime="00:01:16.93" lane="7" heatid="2002" />
                <RESULT resultid="681" eventid="12" swimtime="00:02:44.44" lane="8" heatid="12003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:18.28" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="695" eventid="17" swimtime="00:00:34.95" lane="7" heatid="17002" />
                <RESULT resultid="684" eventid="26" swimtime="00:05:57.77" lane="2" heatid="26002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:20.63" />
                    <SPLIT distance="200" swimtime="00:02:53.24" />
                    <SPLIT distance="300" swimtime="00:04:28.54" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="167" birthdate="1979-01-01" gender="M" lastname="Schubert" firstname="Michael" license="0">
              <RESULTS>
                <RESULT resultid="694" eventid="17" swimtime="00:00:29.27" lane="2" heatid="17004" />
                <RESULT resultid="691" eventid="19" swimtime="00:00:33.35" lane="1" heatid="19003" />
                <RESULT resultid="674" eventid="22" swimtime="00:01:16.56" lane="4" heatid="22001" />
                <RESULT resultid="683" eventid="26" swimtime="00:05:58.67" lane="6" heatid="26002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:16.66" />
                    <SPLIT distance="200" swimtime="00:02:50.35" />
                    <SPLIT distance="300" swimtime="00:04:24.94" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="168" birthdate="1999-01-01" gender="F" lastname="Jacke" firstname="Lena" license="0">
              <RESULTS>
                <RESULT resultid="685" eventid="5" swimtime="00:04:19.93" lane="4" heatid="5001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:59.58" />
                    <SPLIT distance="200" swimtime="00:02:04.50" />
                    <SPLIT distance="300" swimtime="00:03:15.58" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="675" eventid="11" swimtime="00:01:56.54" lane="4" heatid="11009">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:57.73" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="169" birthdate="2005-01-01" gender="M" lastname="Preuß" firstname="Marek" license="0">
              <RESULTS>
                <RESULT resultid="686" eventid="6" swimtime="00:03:36.13" lane="2" heatid="6002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:48.55" />
                    <SPLIT distance="200" swimtime="00:01:44.65" />
                    <SPLIT distance="300" swimtime="00:02:42.31" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="679" eventid="12" swimtime="00:01:45.22" lane="5" heatid="12006">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:52.37" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="SSV Freiburg" nation="GER" region="33" code="0">
          <ATHLETES>
            <ATHLETE athleteid="36" birthdate="1994-01-01" gender="F" lastname="Längin" firstname="Jana" license="0">
              <RESULTS>
                <RESULT resultid="147" eventid="3" swimtime="00:01:04.93" lane="2" heatid="3004" />
                <RESULT resultid="164" eventid="5" swimtime="00:05:06.35" lane="3" heatid="5001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:04.18" />
                    <SPLIT distance="200" swimtime="00:02:21.57" />
                    <SPLIT distance="300" swimtime="00:03:43.64" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="156" eventid="11" swimtime="00:02:24.36" lane="4" heatid="11007">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:08.32" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="170" eventid="16" swimtime="00:00:28.40" lane="1" heatid="16007" />
                <RESULT resultid="168" eventid="18" swimtime="00:00:29.23" lane="2" heatid="18004" />
                <RESULT resultid="152" eventid="21" swimtime="00:00:56.03" lane="4" heatid="21004" />
                <RESULT resultid="160" eventid="25" swimtime="00:05:18.71" lane="7" heatid="25005">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:09.42" />
                    <SPLIT distance="200" swimtime="00:02:31.16" />
                    <SPLIT distance="300" swimtime="00:03:55.82" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="37" birthdate="2000-01-01" gender="F" lastname="Köhn" firstname="Theresa" license="0">
              <RESULTS>
                <RESULT resultid="148" eventid="1" swimtime="00:00:47.49" lane="3" heatid="1012" />
                <RESULT resultid="162" eventid="5" swimtime="00:03:41.88" lane="4" heatid="5002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:52.17" />
                    <SPLIT distance="200" swimtime="00:01:47.54" />
                    <SPLIT distance="300" swimtime="00:02:45.06" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="166" eventid="7" swimtime="00:00:19.78" lane="7" heatid="7005" />
                <RESULT resultid="169" eventid="16" swimtime="00:00:21.59" lane="6" heatid="16011" />
                <RESULT resultid="151" eventid="21" swimtime="00:00:44.46" lane="2" heatid="21006" />
                <RESULT resultid="159" eventid="25" swimtime="00:03:58.93" lane="1" heatid="25008">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:56.83" />
                    <SPLIT distance="200" swimtime="00:01:57.84" />
                    <SPLIT distance="300" swimtime="00:02:59.94" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="38" birthdate="1998-01-01" gender="F" lastname="Köhn" firstname="Johanna" license="0">
              <RESULTS>
                <RESULT resultid="149" eventid="1" swimtime="00:00:47.04" lane="7" heatid="1012" />
                <RESULT resultid="163" eventid="5" swimtime="00:03:45.72" lane="5" heatid="5002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:52.72" />
                    <SPLIT distance="200" swimtime="00:01:49.31" />
                    <SPLIT distance="300" swimtime="00:02:47.74" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="155" eventid="11" swimtime="00:01:43.28" lane="5" heatid="11010">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:50.90" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="154" eventid="15" swimtime="00:15:30.29" lane="5" heatid="15002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:55.55" />
                    <SPLIT distance="200" swimtime="00:01:54.36" />
                    <SPLIT distance="300" swimtime="00:02:54.19" />
                    <SPLIT distance="400" swimtime="00:03:54.87" />
                    <SPLIT distance="500" swimtime="00:04:56.57" />
                    <SPLIT distance="600" swimtime="00:05:59.04" />
                    <SPLIT distance="700" swimtime="00:07:01.88" />
                    <SPLIT distance="800" swimtime="00:08:04.88" />
                    <SPLIT distance="900" swimtime="00:09:08.20" />
                    <SPLIT distance="1000" swimtime="00:10:11.43" />
                    <SPLIT distance="1100" swimtime="00:11:14.74" />
                    <SPLIT distance="1200" swimtime="00:12:18.06" />
                    <SPLIT distance="1300" swimtime="00:13:20.77" />
                    <SPLIT distance="1400" swimtime="00:14:23.06" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="172" eventid="20" swimtime="00:07:58.00" lane="4" heatid="20004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:53.48" />
                    <SPLIT distance="200" swimtime="00:01:51.51" />
                    <SPLIT distance="300" swimtime="00:02:51.91" />
                    <SPLIT distance="400" swimtime="00:03:53.35" />
                    <SPLIT distance="500" swimtime="00:04:55.14" />
                    <SPLIT distance="600" swimtime="00:05:56.99" />
                    <SPLIT distance="700" swimtime="00:06:58.44" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="158" eventid="25" swimtime="00:03:47.13" lane="4" heatid="25008">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:53.56" />
                    <SPLIT distance="200" swimtime="00:01:51.23" />
                    <SPLIT distance="300" swimtime="00:02:49.04" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="39" birthdate="1980-01-01" gender="M" lastname="Schmidt" firstname="Sascha" license="0">
              <RESULTS>
                <RESULT resultid="150" eventid="2" swimtime="00:00:47.32" lane="4" heatid="2007" />
                <RESULT resultid="165" eventid="6" swimtime="00:03:40.19" lane="6" heatid="6002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:50.64" />
                    <SPLIT distance="200" swimtime="00:01:45.00" />
                    <SPLIT distance="300" swimtime="00:02:42.32" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="167" eventid="8" swimtime="00:00:18.62" lane="3" heatid="8003" />
                <RESULT resultid="157" eventid="12" swimtime="00:01:47.26" lane="7" heatid="12007">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:50.75" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="171" eventid="17" swimtime="00:00:21.31" lane="3" heatid="17007" />
                <RESULT resultid="173" eventid="20" swimtime="00:08:41.23" lane="3" heatid="20004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:57.42" />
                    <SPLIT distance="200" swimtime="00:02:01.16" />
                    <SPLIT distance="300" swimtime="00:03:06.54" />
                    <SPLIT distance="400" swimtime="00:04:11.79" />
                    <SPLIT distance="500" swimtime="00:05:18.42" />
                    <SPLIT distance="600" swimtime="00:06:26.03" />
                    <SPLIT distance="700" swimtime="00:07:33.74" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="153" eventid="22" swimtime="00:00:43.27" lane="2" heatid="22004" />
                <RESULT resultid="161" eventid="26" swimtime="00:04:09.23" lane="6" heatid="26005">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:54.83" />
                    <SPLIT distance="200" swimtime="00:01:57.48" />
                    <SPLIT distance="300" swimtime="00:03:03.17" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="Tauchclub Heilbronn" nation="GER" region="32" code="0">
          <ATHLETES>
            <ATHLETE athleteid="40" birthdate="2006-01-01" gender="M" lastname="Cherenok" firstname="Oleksii" license="0">
              <RESULTS>
                <RESULT resultid="174" eventid="4" swimtime="00:00:50.11" lane="5" heatid="4003" />
                <RESULT resultid="248" eventid="8" swimtime="00:00:17.99" lane="5" heatid="8003" />
                <RESULT resultid="252" eventid="19" swimtime="00:00:22.73" lane="5" heatid="19004" />
                <RESULT resultid="201" eventid="22" swimtime="00:00:44.96" lane="8" heatid="22004" />
                <RESULT resultid="226" eventid="26" swimtime="00:04:04.30" lane="2" heatid="26005">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:53.02" />
                    <SPLIT distance="200" swimtime="00:01:54.36" />
                    <SPLIT distance="300" swimtime="00:02:59.42" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="41" birthdate="2004-01-01" gender="F" lastname="Phillipp" firstname="Beeke Alea" license="0">
              <RESULTS>
                <RESULT resultid="175" eventid="1" swimtime="00:00:47.73" lane="6" heatid="1012" />
                <RESULT resultid="240" eventid="7" swimtime="00:00:19.84" lane="5" heatid="7004" />
                <RESULT resultid="258" eventid="16" swimtime="00:00:21.27" lane="7" heatid="16011" />
                <RESULT resultid="193" eventid="21" swimtime="00:00:45.53" lane="4" heatid="21005" />
                <RESULT resultid="216" eventid="25" swimtime="00:03:58.38" lane="8" heatid="25008">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:53.01" />
                    <SPLIT distance="200" swimtime="00:01:51.93" />
                    <SPLIT distance="300" swimtime="00:02:55.63" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="42" birthdate="2009-01-01" gender="F" lastname="Hölzer" firstname="Elisa" license="0">
              <RESULTS>
                <RESULT resultid="176" eventid="1" swimtime="00:00:52.59" lane="5" heatid="1010" />
                <RESULT resultid="241" eventid="7" swimtime="00:00:21.57" lane="6" heatid="7003" />
                <RESULT resultid="205" eventid="11" swimtime="00:01:56.18" lane="2" heatid="11009">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:54.46" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="260" eventid="16" swimtime="00:00:23.66" lane="2" heatid="16010" />
                <RESULT resultid="195" eventid="21" swimtime="00:00:53.52" lane="7" heatid="21005" />
                <RESULT resultid="218" eventid="25" swimtime="00:04:17.15" lane="2" heatid="25007">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:58.42" />
                    <SPLIT distance="200" swimtime="00:02:05.80" />
                    <SPLIT distance="300" swimtime="00:03:13.78" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="43" birthdate="2000-01-01" gender="F" lastname="Baier" firstname="Jessika" license="0">
              <RESULTS>
                <RESULT resultid="177" eventid="1" swimtime="00:00:54.78" lane="6" heatid="1010" />
                <RESULT resultid="244" eventid="7" swimtime="00:00:21.56" lane="8" heatid="7003" />
                <RESULT resultid="263" eventid="16" swimtime="00:00:23.82" lane="2" heatid="16009" />
                <RESULT resultid="196" eventid="21" swimtime="00:00:52.12" lane="5" heatid="21004" />
                <RESULT resultid="219" eventid="25" swimtime="00:04:40.54" lane="4" heatid="25006">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:56.59" />
                    <SPLIT distance="200" swimtime="00:02:08.03" />
                    <SPLIT distance="300" swimtime="00:03:25.22" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="44" birthdate="2008-01-01" gender="F" lastname="Seidel" firstname="Esther-Sophie" license="0">
              <RESULTS>
                <RESULT resultid="178" eventid="1" swimtime="00:00:52.14" lane="2" heatid="1010" />
                <RESULT resultid="242" eventid="7" swimtime="00:00:21.10" lane="2" heatid="7003" />
                <RESULT resultid="261" eventid="16" swimtime="00:00:22.48" lane="1" heatid="16010" />
                <RESULT resultid="198" eventid="21" swimtime="00:00:56.89" lane="4" heatid="21003" />
                <RESULT resultid="220" eventid="25" status="DSQ" swimtime="00:04:26.11" lane="5" heatid="25006" comment="falscher Start">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:57.68" />
                    <SPLIT distance="200" swimtime="00:02:09.17" />
                    <SPLIT distance="300" swimtime="00:03:19.89" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="45" birthdate="2008-01-01" gender="F" lastname="Grimm" firstname="Hannah" license="0">
              <RESULTS>
                <RESULT resultid="179" eventid="1" status="DNS" swimtime="00:00:00.00" lane="8" heatid="1009" />
                <RESULT resultid="243" eventid="7" status="DNS" swimtime="00:00:00.00" lane="7" heatid="7003" />
                <RESULT resultid="262" eventid="16" status="DNS" swimtime="00:00:00.00" lane="8" heatid="16010" />
                <RESULT resultid="197" eventid="21" status="DNS" swimtime="00:00:00.00" lane="1" heatid="21004" />
                <RESULT resultid="221" eventid="25" status="DNS" swimtime="00:00:00.00" lane="6" heatid="25006" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="46" birthdate="2009-01-01" gender="F" lastname="Rettig" firstname="Sina" license="0">
              <RESULTS>
                <RESULT resultid="180" eventid="1" swimtime="00:00:58.32" lane="3" heatid="1008" />
                <RESULT resultid="245" eventid="7" swimtime="00:00:24.59" lane="5" heatid="7002" />
                <RESULT resultid="206" eventid="11" swimtime="00:02:16.18" lane="5" heatid="11007">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:05.22" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="264" eventid="16" swimtime="00:00:25.43" lane="6" heatid="16008" />
                <RESULT resultid="199" eventid="21" swimtime="00:01:02.44" lane="7" heatid="21003" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="47" birthdate="2012-01-01" gender="F" lastname="Grimmig" firstname="Jella" license="0">
              <RESULTS>
                <RESULT resultid="181" eventid="1" swimtime="00:01:02.36" lane="8" heatid="1007" />
                <RESULT resultid="208" eventid="11" swimtime="00:02:24.95" lane="2" heatid="11006">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:09.93" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="266" eventid="16" swimtime="00:00:27.59" lane="6" heatid="16005" />
                <RESULT resultid="254" eventid="23" swimtime="00:00:30.30" lane="3" heatid="23004" />
                <RESULT resultid="222" eventid="25" swimtime="00:05:08.57" lane="5" heatid="25004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:08.38" />
                    <SPLIT distance="200" swimtime="00:02:29.65" />
                    <SPLIT distance="300" swimtime="00:03:51.59" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="48" birthdate="2012-01-01" gender="F" lastname="Leleux" firstname="Frida Julie" license="0">
              <RESULTS>
                <RESULT resultid="182" eventid="1" swimtime="00:01:00.73" lane="1" heatid="1006" />
                <RESULT resultid="207" eventid="11" swimtime="00:02:21.72" lane="6" heatid="11006">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:05.84" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="265" eventid="16" status="DSQ" swimtime="00:00:26.95" lane="7" heatid="16006" comment="falscher Start" />
                <RESULT resultid="253" eventid="23" swimtime="00:00:31.79" lane="5" heatid="23004" />
                <RESULT resultid="224" eventid="25" swimtime="00:05:24.82" lane="5" heatid="25003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:06.98" />
                    <SPLIT distance="200" swimtime="00:02:31.24" />
                    <SPLIT distance="300" swimtime="00:04:00.81" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="49" birthdate="2011-01-01" gender="F" lastname="Jung" firstname="Sarah" license="0">
              <RESULTS>
                <RESULT resultid="183" eventid="1" swimtime="00:01:06.93" lane="5" heatid="1005" />
                <RESULT resultid="209" eventid="11" swimtime="00:02:31.02" lane="6" heatid="11005">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:14.05" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="267" eventid="16" swimtime="00:00:29.58" lane="7" heatid="16005" />
                <RESULT resultid="223" eventid="25" swimtime="00:05:35.37" lane="2" heatid="25004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:15.68" />
                    <SPLIT distance="200" swimtime="00:02:45.15" />
                    <SPLIT distance="300" swimtime="00:04:09.72" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="50" birthdate="2014-01-01" gender="F" lastname="Nagel" firstname="Marlene" license="0">
              <RESULTS>
                <RESULT resultid="184" eventid="1" swimtime="00:01:36.09" lane="4" heatid="1001" />
                <RESULT resultid="210" eventid="11" swimtime="00:03:34.83" lane="8" heatid="11002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:42.88" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="268" eventid="16" swimtime="00:00:38.56" lane="5" heatid="16001" />
                <RESULT resultid="251" eventid="18" swimtime="00:00:40.90" lane="7" heatid="18002" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="51" birthdate="2003-01-01" gender="M" lastname="Fabriz" firstname="Tobias" license="0">
              <RESULTS>
                <RESULT resultid="185" eventid="2" swimtime="00:00:43.41" lane="1" heatid="2008" />
                <RESULT resultid="246" eventid="8" swimtime="00:00:17.06" lane="7" heatid="8004" />
                <RESULT resultid="269" eventid="17" swimtime="00:00:19.21" lane="8" heatid="17008" />
                <RESULT resultid="200" eventid="22" swimtime="00:00:41.63" lane="6" heatid="22004" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="54" birthdate="2002-01-01" gender="M" lastname="Bauer" firstname="Sebastian" license="0">
              <RESULTS>
                <RESULT resultid="188" eventid="2" swimtime="00:00:51.81" lane="7" heatid="2006" />
                <RESULT resultid="249" eventid="8" swimtime="00:00:19.75" lane="5" heatid="8002" />
                <RESULT resultid="212" eventid="12" swimtime="00:01:56.93" lane="2" heatid="12006">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:56.43" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="272" eventid="17" swimtime="00:00:22.89" lane="5" heatid="17006" />
                <RESULT resultid="228" eventid="26" swimtime="00:04:12.45" lane="4" heatid="26004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:57.63" />
                    <SPLIT distance="200" swimtime="00:02:01.56" />
                    <SPLIT distance="300" swimtime="00:03:07.85" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="55" birthdate="2011-01-01" gender="M" lastname="Korb" firstname="Elias" license="0">
              <RESULTS>
                <RESULT resultid="189" eventid="2" swimtime="00:00:58.40" lane="7" heatid="2005" />
                <RESULT resultid="277" eventid="10" swimtime="00:00:24.64" lane="5" heatid="10002" />
                <RESULT resultid="273" eventid="17" swimtime="00:00:26.34" lane="4" heatid="17004" />
                <RESULT resultid="203" eventid="22" swimtime="00:00:56.24" lane="3" heatid="22002" />
                <RESULT resultid="229" eventid="26" swimtime="00:04:21.10" lane="3" heatid="26004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:02.55" />
                    <SPLIT distance="200" swimtime="00:02:10.16" />
                    <SPLIT distance="300" swimtime="00:03:18.97" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="56" birthdate="2012-01-01" gender="M" lastname="Hölzer" firstname="Vincent" license="0">
              <RESULTS>
                <RESULT resultid="190" eventid="2" swimtime="00:01:06.53" lane="8" heatid="2004" />
                <RESULT resultid="213" eventid="12" swimtime="00:02:28.77" lane="1" heatid="12004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:12.49" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="274" eventid="17" swimtime="00:00:30.32" lane="7" heatid="17004" />
                <RESULT resultid="255" eventid="24" swimtime="00:00:33.22" lane="4" heatid="24002" />
                <RESULT resultid="230" eventid="26" swimtime="00:05:14.71" lane="8" heatid="26003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:13.60" />
                    <SPLIT distance="200" swimtime="00:02:37.16" />
                    <SPLIT distance="300" swimtime="00:03:56.55" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="57" birthdate="2013-01-01" gender="M" lastname="Lang" firstname="Leo" license="0">
              <RESULTS>
                <RESULT resultid="191" eventid="2" swimtime="00:01:11.04" lane="5" heatid="2002" />
                <RESULT resultid="214" eventid="12" swimtime="00:02:42.43" lane="2" heatid="12003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:15.87" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="276" eventid="17" swimtime="00:00:29.94" lane="4" heatid="17002" />
                <RESULT resultid="257" eventid="24" swimtime="00:00:35.76" lane="2" heatid="24002" />
                <RESULT resultid="231" eventid="26" swimtime="00:05:59.20" lane="8" heatid="26002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:23.85" />
                    <SPLIT distance="200" swimtime="00:03:02.57" />
                    <SPLIT distance="300" swimtime="00:04:37.75" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="58" birthdate="2013-01-01" gender="M" lastname="Phillipp" firstname="Daan Iven" license="0">
              <RESULTS>
                <RESULT resultid="192" eventid="2" swimtime="00:01:21.49" lane="6" heatid="2002" />
                <RESULT resultid="215" eventid="12" swimtime="00:02:46.41" lane="5" heatid="12002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:18.08" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="275" eventid="17" swimtime="00:00:33.77" lane="8" heatid="17003" />
                <RESULT resultid="256" eventid="24" swimtime="00:00:38.08" lane="6" heatid="24002" />
                <RESULT resultid="232" eventid="26" swimtime="00:06:28.01" lane="4" heatid="26001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:26.74" />
                    <SPLIT distance="200" swimtime="00:03:07.89" />
                    <SPLIT distance="300" swimtime="00:04:48.96" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="59" birthdate="2004-01-01" gender="F" lastname="Ruedel" firstname="Leona" license="0">
              <RESULTS>
                <RESULT resultid="239" eventid="7" swimtime="00:00:19.27" lane="8" heatid="7005" />
                <RESULT resultid="204" eventid="11" swimtime="00:01:46.96" lane="6" heatid="11010">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:51.68" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="259" eventid="16" swimtime="00:00:21.80" lane="5" heatid="16010" />
                <RESULT resultid="194" eventid="21" swimtime="00:00:45.83" lane="3" heatid="21005" />
                <RESULT resultid="217" eventid="25" swimtime="00:03:55.60" lane="4" heatid="25007">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:53.32" />
                    <SPLIT distance="200" swimtime="00:01:54.07" />
                    <SPLIT distance="300" swimtime="00:02:56.79" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY number="1" gender="F" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="233" eventid="28" swimtime="00:03:49.26" lane="6" heatid="28001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:53.60" />
                    <SPLIT distance="200" swimtime="00:01:57.29" />
                    <SPLIT distance="300" swimtime="00:02:58.54" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="42" number="1" />
                    <RELAYPOSITION athleteid="48" number="2" />
                    <RELAYPOSITION athleteid="46" number="3" />
                    <RELAYPOSITION athleteid="44" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" gender="M" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="235" eventid="29" swimtime="00:04:37.12" lane="1" heatid="29001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:06.96" />
                    <SPLIT distance="200" swimtime="00:02:19.06" />
                    <SPLIT distance="300" swimtime="00:03:39.12" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="56" number="1" />
                    <RELAYPOSITION athleteid="57" number="2" />
                    <RELAYPOSITION athleteid="58" number="3" />
                    <RELAYPOSITION athleteid="55" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" gender="X" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="237" eventid="13" swimtime="00:01:31.64" lane="7" heatid="13003">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="44" number="1" />
                    <RELAYPOSITION athleteid="55" number="2" />
                    <RELAYPOSITION athleteid="42" number="3" />
                    <RELAYPOSITION athleteid="40" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" gender="X" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="238" eventid="13" swimtime="00:01:55.50" lane="2" heatid="13002">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="47" number="1" />
                    <RELAYPOSITION athleteid="56" number="2" />
                    <RELAYPOSITION athleteid="48" number="3" />
                    <RELAYPOSITION athleteid="57" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB name="Tauchsportclub Erfurt e.V." nation="GER" region="35" code="0">
          <ATHLETES>
            <ATHLETE athleteid="184" birthdate="2009-01-01" gender="F" lastname="Blumenstein" firstname="Martha" license="0">
              <RESULTS>
                <RESULT resultid="768" eventid="3" swimtime="00:00:57.94" lane="4" heatid="3004" />
                <RESULT resultid="884" eventid="7" swimtime="00:00:23.63" lane="5" heatid="7001" />
                <RESULT resultid="823" eventid="11" swimtime="00:02:09.00" lane="2" heatid="11008">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:02.68" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="818" eventid="15" swimtime="00:18:52.40" lane="4" heatid="15001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:06.32" />
                    <SPLIT distance="200" swimtime="00:02:21.27" />
                    <SPLIT distance="300" swimtime="00:03:37.06" />
                    <SPLIT distance="400" swimtime="00:04:53.61" />
                    <SPLIT distance="500" swimtime="00:06:11.96" />
                    <SPLIT distance="600" swimtime="00:07:27.91" />
                    <SPLIT distance="700" swimtime="00:08:45.36" />
                    <SPLIT distance="800" swimtime="00:10:02.32" />
                    <SPLIT distance="900" swimtime="00:11:19.84" />
                    <SPLIT distance="1000" swimtime="00:12:36.41" />
                    <SPLIT distance="1100" swimtime="00:13:53.47" />
                    <SPLIT distance="1200" swimtime="00:15:10.95" />
                    <SPLIT distance="1300" swimtime="00:16:26.94" />
                    <SPLIT distance="1400" swimtime="00:17:41.77" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="921" eventid="16" swimtime="00:00:24.15" lane="8" heatid="16008" />
                <RESULT resultid="892" eventid="18" swimtime="00:00:26.75" lane="7" heatid="18005" />
                <RESULT resultid="950" eventid="20" swimtime="00:09:58.10" lane="8" heatid="20003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:07.12" />
                    <SPLIT distance="200" swimtime="00:02:22.32" />
                    <SPLIT distance="300" swimtime="00:03:37.67" />
                    <SPLIT distance="400" swimtime="00:04:53.27" />
                    <SPLIT distance="500" swimtime="00:06:08.06" />
                    <SPLIT distance="600" swimtime="00:07:24.55" />
                    <SPLIT distance="700" swimtime="00:08:41.69" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="185" birthdate="1982-01-01" gender="F" lastname="Zitzmann" firstname="Ulrike" license="0">
              <RESULTS>
                <RESULT resultid="789" eventid="1" swimtime="00:01:07.18" lane="3" heatid="1007" />
                <RESULT resultid="769" eventid="3" swimtime="00:01:07.46" lane="5" heatid="3004" />
                <RESULT resultid="925" eventid="16" swimtime="00:00:27.96" lane="4" heatid="16006" />
                <RESULT resultid="893" eventid="18" swimtime="00:00:27.79" lane="1" heatid="18005" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="186" birthdate="2009-01-01" gender="F" lastname="Henkel" firstname="Friederike" license="0">
              <RESULTS>
                <RESULT resultid="792" eventid="1" swimtime="00:01:01.45" lane="3" heatid="1006" />
                <RESULT resultid="770" eventid="3" swimtime="00:01:09.84" lane="7" heatid="3004" />
                <RESULT resultid="826" eventid="11" swimtime="00:02:19.86" lane="4" heatid="11006">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:06.21" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="923" eventid="16" swimtime="00:00:25.84" lane="2" heatid="16007" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="187" birthdate="2007-01-01" gender="F" lastname="Zieger" firstname="Emilie" license="0">
              <RESULTS>
                <RESULT resultid="790" eventid="1" status="DNS" swimtime="00:00:00.00" lane="6" heatid="1007" />
                <RESULT resultid="771" eventid="3" status="DNS" swimtime="00:00:00.00" lane="4" heatid="3003" />
                <RESULT resultid="825" eventid="11" status="DNS" swimtime="00:00:00.00" lane="2" heatid="11007" />
                <RESULT resultid="926" eventid="16" swimtime="00:00:28.73" lane="8" heatid="16006" />
                <RESULT resultid="850" eventid="25" status="DSQ" swimtime="00:00:00.00" lane="8" heatid="25005" comment="aufgegeben nach 140m">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:09.06" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="188" birthdate="2012-01-01" gender="F" lastname="Palchyk" firstname="Myroslava" license="0">
              <RESULTS>
                <RESULT resultid="794" eventid="1" swimtime="00:01:06.70" lane="1" heatid="1005" />
                <RESULT resultid="772" eventid="3" swimtime="00:01:08.89" lane="5" heatid="3003" />
                <RESULT resultid="829" eventid="11" swimtime="00:02:35.29" lane="3" heatid="11005">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:12.04" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="932" eventid="16" swimtime="00:00:28.89" lane="3" heatid="16002" />
                <RESULT resultid="897" eventid="18" swimtime="00:00:30.59" lane="2" heatid="18003" />
                <RESULT resultid="909" eventid="23" swimtime="00:00:30.39" lane="2" heatid="23004" />
                <RESULT resultid="854" eventid="25" swimtime="00:05:40.37" lane="3" heatid="25003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:17.74" />
                    <SPLIT distance="200" swimtime="00:02:51.19" />
                    <SPLIT distance="300" swimtime="00:04:13.51" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="189" birthdate="2012-01-01" gender="F" lastname="Blumenstein" firstname="Liese" license="0">
              <RESULTS>
                <RESULT resultid="793" eventid="1" swimtime="00:01:15.45" lane="2" heatid="1005" />
                <RESULT resultid="773" eventid="3" swimtime="00:01:12.13" lane="3" heatid="3003" />
                <RESULT resultid="828" eventid="11" swimtime="00:02:34.81" lane="4" heatid="11005">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:16.37" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="931" eventid="16" swimtime="00:00:32.44" lane="1" heatid="16003" />
                <RESULT resultid="896" eventid="18" swimtime="00:00:30.62" lane="8" heatid="18004" />
                <RESULT resultid="908" eventid="23" swimtime="00:00:34.02" lane="6" heatid="23004" />
                <RESULT resultid="853" eventid="25" swimtime="00:05:33.75" lane="8" heatid="25004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:18.41" />
                    <SPLIT distance="200" swimtime="00:02:47.22" />
                    <SPLIT distance="300" swimtime="00:04:13.87" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="190" birthdate="2011-01-01" gender="F" lastname="Döll" firstname="Katharina Martha" license="0">
              <RESULTS>
                <RESULT resultid="796" eventid="1" status="DSQ" swimtime="00:00:00.00" lane="4" heatid="1003" comment="Aufgegeben nach 50 m" />
                <RESULT resultid="774" eventid="3" swimtime="00:01:13.25" lane="1" heatid="3003" />
                <RESULT resultid="831" eventid="11" swimtime="00:02:40.84" lane="8" heatid="11003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:17.72" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="929" eventid="16" swimtime="00:00:36.41" lane="2" heatid="16003" />
                <RESULT resultid="855" eventid="25" swimtime="00:05:37.32" lane="1" heatid="25003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:15.17" />
                    <SPLIT distance="200" swimtime="00:02:44.72" />
                    <SPLIT distance="300" swimtime="00:04:13.55" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="191" birthdate="2013-01-01" gender="F" lastname="Medola" firstname="Anna" license="0">
              <RESULTS>
                <RESULT resultid="775" eventid="3" swimtime="00:01:31.62" lane="7" heatid="3002" />
                <RESULT resultid="833" eventid="11" swimtime="00:03:28.60" lane="1" heatid="11002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:43.30" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="899" eventid="18" swimtime="00:00:36.56" lane="6" heatid="18002" />
                <RESULT resultid="912" eventid="23" swimtime="00:00:44.59" lane="6" heatid="23002" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="192" birthdate="2013-01-01" gender="F" lastname="Hohmann" firstname="Jette" license="0">
              <RESULTS>
                <RESULT resultid="776" eventid="3" swimtime="00:01:23.63" lane="1" heatid="3002" />
                <RESULT resultid="834" eventid="11" swimtime="00:03:20.10" lane="5" heatid="11001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:42.58" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="898" eventid="18" swimtime="00:00:35.85" lane="3" heatid="18002" />
                <RESULT resultid="907" eventid="23" swimtime="00:00:38.94" lane="3" heatid="23001" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="194" birthdate="2009-01-01" gender="M" lastname="Artschwager" firstname="Gustaf" license="0">
              <RESULTS>
                <RESULT resultid="778" eventid="4" swimtime="00:00:58.85" lane="4" heatid="4002" />
                <RESULT resultid="839" eventid="12" swimtime="00:02:11.54" lane="1" heatid="12005">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:03.79" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="817" eventid="15" swimtime="00:20:26.45" lane="6" heatid="15001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:12.11" />
                    <SPLIT distance="200" swimtime="00:02:33.92" />
                    <SPLIT distance="300" swimtime="00:03:56.55" />
                    <SPLIT distance="400" swimtime="00:05:18.59" />
                    <SPLIT distance="500" swimtime="00:06:42.50" />
                    <SPLIT distance="600" swimtime="00:08:06.56" />
                    <SPLIT distance="700" swimtime="00:09:30.36" />
                    <SPLIT distance="800" swimtime="00:10:54.70" />
                    <SPLIT distance="900" swimtime="00:12:19.57" />
                    <SPLIT distance="1000" swimtime="00:13:42.50" />
                    <SPLIT distance="1100" swimtime="00:15:06.10" />
                    <SPLIT distance="1200" swimtime="00:16:29.42" />
                    <SPLIT distance="1300" swimtime="00:17:52.59" />
                    <SPLIT distance="1400" swimtime="00:19:12.36" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="940" eventid="17" swimtime="00:00:28.19" lane="5" heatid="17004" />
                <RESULT resultid="951" eventid="20" swimtime="00:10:18.55" lane="5" heatid="20002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:05.00" />
                    <SPLIT distance="200" swimtime="00:02:21.87" />
                    <SPLIT distance="300" swimtime="00:03:41.23" />
                    <SPLIT distance="400" swimtime="00:05:00.54" />
                    <SPLIT distance="500" swimtime="00:06:21.31" />
                    <SPLIT distance="600" swimtime="00:07:42.57" />
                    <SPLIT distance="700" swimtime="00:09:02.65" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="816" eventid="22" swimtime="00:01:09.44" lane="6" heatid="22001" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="195" birthdate="2010-01-01" gender="M" lastname="Schmidt" firstname="Jakob" license="0">
              <RESULTS>
                <RESULT resultid="779" eventid="4" swimtime="00:01:12.97" lane="1" heatid="4002" />
                <RESULT resultid="843" eventid="12" swimtime="00:02:47.15" lane="6" heatid="12003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:20.60" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="942" eventid="17" swimtime="00:00:32.71" lane="2" heatid="17003" />
                <RESULT resultid="903" eventid="19" swimtime="00:00:30.63" lane="3" heatid="19002" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="196" birthdate="2012-01-01" gender="M" lastname="Geyer" firstname="Julius" license="0">
              <RESULTS>
                <RESULT resultid="807" eventid="2" swimtime="00:01:22.03" lane="4" heatid="2002" />
                <RESULT resultid="780" eventid="4" swimtime="00:01:23.85" lane="8" heatid="4002" />
                <RESULT resultid="845" eventid="12" swimtime="00:03:02.94" lane="2" heatid="12002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:28.06" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="943" eventid="17" swimtime="00:00:36.60" lane="6" heatid="17002" />
                <RESULT resultid="906" eventid="19" swimtime="00:00:37.60" lane="2" heatid="19001" />
                <RESULT resultid="913" eventid="24" swimtime="00:00:39.12" lane="3" heatid="24002" />
                <RESULT resultid="859" eventid="26" swimtime="00:06:34.14" lane="2" heatid="26001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:27.85" />
                    <SPLIT distance="200" swimtime="00:03:08.13" />
                    <SPLIT distance="300" swimtime="00:04:55.52" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="197" birthdate="2014-01-01" gender="M" lastname="Schmidt" firstname="Arthur" license="0">
              <RESULTS>
                <RESULT resultid="781" eventid="4" swimtime="00:01:21.68" lane="5" heatid="4001" />
                <RESULT resultid="844" eventid="12" swimtime="00:02:58.42" lane="6" heatid="12002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:26.24" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="904" eventid="19" swimtime="00:00:37.00" lane="5" heatid="19001" />
                <RESULT resultid="914" eventid="24" swimtime="00:00:42.37" lane="3" heatid="24001" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="198" birthdate="2011-01-01" gender="M" lastname="Heidrich" firstname="Pascal" license="0">
              <RESULTS>
                <RESULT resultid="782" eventid="4" swimtime="00:01:34.82" lane="7" heatid="4001" />
                <RESULT resultid="835" eventid="12" status="DSQ" swimtime="00:04:15.96" lane="3" heatid="12001" comment="falsche Schwimmtechnik (keine Schnorchelatmung, Regelwerk CMAS 2.2.1.4)">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:44.30" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="905" eventid="19" status="DNS" swimtime="00:00:00.00" lane="3" heatid="19001" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="199" birthdate="2009-01-01" gender="F" lastname="Darzhaniia" firstname="Alisa" license="0">
              <RESULTS>
                <RESULT resultid="783" eventid="1" swimtime="00:00:48.41" lane="5" heatid="1011" />
                <RESULT resultid="879" eventid="7" swimtime="00:00:19.90" lane="3" heatid="7004" />
                <RESULT resultid="820" eventid="11" swimtime="00:01:49.71" lane="1" heatid="11010">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:52.26" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="915" eventid="16" swimtime="00:00:22.13" lane="8" heatid="16011" />
                <RESULT resultid="890" eventid="18" swimtime="00:00:25.58" lane="4" heatid="18005" />
                <RESULT resultid="949" eventid="20" swimtime="00:08:22.09" lane="7" heatid="20004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:56.03" />
                    <SPLIT distance="200" swimtime="00:01:59.02" />
                    <SPLIT distance="300" swimtime="00:03:03.63" />
                    <SPLIT distance="400" swimtime="00:04:08.52" />
                    <SPLIT distance="500" swimtime="00:05:13.75" />
                    <SPLIT distance="600" swimtime="00:06:18.70" />
                    <SPLIT distance="700" swimtime="00:07:22.14" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="201" birthdate="2006-01-01" gender="F" lastname="Heinitz" firstname="Leonor" license="0">
              <RESULTS>
                <RESULT resultid="785" eventid="1" swimtime="00:00:53.99" lane="7" heatid="1010" />
                <RESULT resultid="881" eventid="7" swimtime="00:00:21.71" lane="5" heatid="7003" />
                <RESULT resultid="821" eventid="11" swimtime="00:02:01.53" lane="6" heatid="11009">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:57.11" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="917" eventid="16" swimtime="00:00:24.04" lane="4" heatid="16009" />
                <RESULT resultid="808" eventid="21" swimtime="00:00:51.63" lane="1" heatid="21005" />
                <RESULT resultid="846" eventid="25" swimtime="00:04:19.77" lane="3" heatid="25007">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:58.02" />
                    <SPLIT distance="200" swimtime="00:02:05.46" />
                    <SPLIT distance="300" swimtime="00:03:14.27" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="202" birthdate="2010-01-01" gender="F" lastname="Abe" firstname="Adina" license="0">
              <RESULTS>
                <RESULT resultid="786" eventid="1" swimtime="00:00:51.60" lane="8" heatid="1010" />
                <RESULT resultid="945" eventid="9" swimtime="00:00:23.62" lane="4" heatid="9002" />
                <RESULT resultid="822" eventid="11" swimtime="00:01:58.56" lane="7" heatid="11009">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:57.59" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="918" eventid="16" swimtime="00:00:23.49" lane="5" heatid="16009" />
                <RESULT resultid="810" eventid="21" swimtime="00:00:50.66" lane="2" heatid="21004" />
                <RESULT resultid="847" eventid="25" swimtime="00:04:18.21" lane="1" heatid="25007">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:00.43" />
                    <SPLIT distance="200" swimtime="00:02:09.04" />
                    <SPLIT distance="300" swimtime="00:03:15.67" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="203" birthdate="2004-01-01" gender="F" lastname="Möller" firstname="Amelie" license="0">
              <RESULTS>
                <RESULT resultid="787" eventid="1" swimtime="00:00:57.44" lane="6" heatid="1009" />
                <RESULT resultid="882" eventid="7" swimtime="00:00:24.82" lane="8" heatid="7002" />
                <RESULT resultid="920" eventid="16" status="DSQ" swimtime="00:00:25.33" lane="4" heatid="16008" comment="falscher Start" />
                <RESULT resultid="894" eventid="18" swimtime="00:00:28.96" lane="5" heatid="18004" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="204" birthdate="1979-01-01" gender="F" lastname="Leipold" firstname="Steffi" license="0">
              <RESULTS>
                <RESULT resultid="788" eventid="1" swimtime="00:00:58.01" lane="2" heatid="1008" />
                <RESULT resultid="883" eventid="7" swimtime="00:00:26.23" lane="4" heatid="7001" />
                <RESULT resultid="824" eventid="11" swimtime="00:02:10.05" lane="7" heatid="11008">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:01.01" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="922" eventid="16" swimtime="00:00:27.01" lane="4" heatid="16007" />
                <RESULT resultid="848" eventid="25" swimtime="00:04:42.78" lane="2" heatid="25006">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:01.97" />
                    <SPLIT distance="200" swimtime="00:02:15.70" />
                    <SPLIT distance="300" swimtime="00:03:30.76" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="205" birthdate="2011-01-01" gender="F" lastname="Behrmann" firstname="Fine Erna" license="0">
              <RESULTS>
                <RESULT resultid="791" eventid="1" swimtime="00:01:04.22" lane="5" heatid="1006" />
                <RESULT resultid="944" eventid="9" swimtime="00:00:30.63" lane="3" heatid="9001" />
                <RESULT resultid="827" eventid="11" swimtime="00:02:27.91" lane="7" heatid="11006">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:08.58" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="924" eventid="16" swimtime="00:00:29.49" lane="8" heatid="16007" />
                <RESULT resultid="852" eventid="25" swimtime="00:05:13.96" lane="1" heatid="25004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:10.95" />
                    <SPLIT distance="200" swimtime="00:02:34.21" />
                    <SPLIT distance="300" swimtime="00:03:58.92" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="206" birthdate="2012-01-01" gender="F" lastname="Schulze" firstname="Paula" license="0">
              <RESULTS>
                <RESULT resultid="795" eventid="1" swimtime="00:01:15.12" lane="6" heatid="1004" />
                <RESULT resultid="830" eventid="11" swimtime="00:02:47.15" lane="5" heatid="11003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:19.09" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="928" eventid="16" swimtime="00:00:32.69" lane="7" heatid="16004" />
                <RESULT resultid="910" eventid="23" swimtime="00:00:34.99" lane="7" heatid="23004" />
                <RESULT resultid="856" eventid="25" swimtime="00:06:04.91" lane="5" heatid="25002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:24.20" />
                    <SPLIT distance="200" swimtime="00:03:01.46" />
                    <SPLIT distance="300" swimtime="00:04:38.85" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="207" birthdate="2010-01-01" gender="F" lastname="Hartung" firstname="Antonia Lea" license="0">
              <RESULTS>
                <RESULT resultid="797" eventid="1" swimtime="00:01:20.61" lane="1" heatid="1003" />
                <RESULT resultid="819" eventid="11" swimtime="00:02:52.07" lane="7" heatid="11001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:22.60" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="930" eventid="16" swimtime="00:00:34.17" lane="7" heatid="16003" />
                <RESULT resultid="857" eventid="25" swimtime="00:06:30.75" lane="4" heatid="25001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:27.63" />
                    <SPLIT distance="200" swimtime="00:03:09.10" />
                    <SPLIT distance="300" swimtime="00:04:49.03" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="208" birthdate="2012-01-01" gender="F" lastname="Dallgas" firstname="Tia" license="0">
              <RESULTS>
                <RESULT resultid="798" eventid="1" swimtime="00:01:10.39" lane="4" heatid="1002" />
                <RESULT resultid="832" eventid="11" swimtime="00:02:43.64" lane="3" heatid="11002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:22.61" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="927" eventid="16" swimtime="00:00:31.47" lane="3" heatid="16004" />
                <RESULT resultid="911" eventid="23" swimtime="00:00:37.88" lane="8" heatid="23004" />
                <RESULT resultid="858" eventid="25" swimtime="00:05:46.93" lane="5" heatid="25001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:25.90" />
                    <SPLIT distance="200" swimtime="00:02:55.47" />
                    <SPLIT distance="300" swimtime="00:04:26.50" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="209" birthdate="2006-01-01" gender="M" lastname="Leipold" firstname="Marek" license="0">
              <RESULTS>
                <RESULT resultid="799" eventid="2" swimtime="00:00:36.46" lane="5" heatid="2008" />
                <RESULT resultid="885" eventid="8" swimtime="00:00:15.53" lane="5" heatid="8004" />
                <RESULT resultid="836" eventid="12" swimtime="00:01:30.87" lane="5" heatid="12007">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:43.29" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="933" eventid="17" swimtime="00:00:16.67" lane="4" heatid="17008" />
                <RESULT resultid="811" eventid="22" swimtime="00:00:35.90" lane="4" heatid="22004" />
                <RESULT resultid="860" eventid="26" swimtime="00:03:20.86" lane="4" heatid="26005">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:45.46" />
                    <SPLIT distance="200" swimtime="00:01:37.53" />
                    <SPLIT distance="300" swimtime="00:02:30.86" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="210" birthdate="1970-01-01" gender="M" lastname="Timpel" firstname="Heiko" license="0">
              <RESULTS>
                <RESULT resultid="800" eventid="2" swimtime="00:00:50.37" lane="1" heatid="2007" />
                <RESULT resultid="866" eventid="6" swimtime="00:03:56.09" lane="1" heatid="6002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:50.00" />
                    <SPLIT distance="200" swimtime="00:01:49.29" />
                    <SPLIT distance="300" swimtime="00:02:53.00" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="886" eventid="8" swimtime="00:00:20.90" lane="8" heatid="8003" />
                <RESULT resultid="934" eventid="17" swimtime="00:00:23.41" lane="4" heatid="17006" />
                <RESULT resultid="900" eventid="19" swimtime="00:00:25.51" lane="5" heatid="19003" />
                <RESULT resultid="812" eventid="22" swimtime="00:00:45.33" lane="4" heatid="22003" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="211" birthdate="2008-01-01" gender="M" lastname="Hannemann" firstname="Fynn" license="0">
              <RESULTS>
                <RESULT resultid="801" eventid="2" swimtime="00:00:50.28" lane="2" heatid="2006" />
                <RESULT resultid="887" eventid="8" swimtime="00:00:22.21" lane="3" heatid="8002" />
                <RESULT resultid="838" eventid="12" swimtime="00:01:59.79" lane="3" heatid="12005">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:57.21" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="935" eventid="17" swimtime="00:00:22.84" lane="6" heatid="17006" />
                <RESULT resultid="814" eventid="22" swimtime="00:00:53.17" lane="4" heatid="22002" />
                <RESULT resultid="862" eventid="26" swimtime="00:04:31.12" lane="8" heatid="26004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:03.80" />
                    <SPLIT distance="200" swimtime="00:02:15.01" />
                    <SPLIT distance="300" swimtime="00:03:26.66" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="212" birthdate="2010-01-01" gender="M" lastname="Leipold" firstname="Jakob" license="0">
              <RESULTS>
                <RESULT resultid="802" eventid="2" swimtime="00:00:55.48" lane="8" heatid="2006" />
                <RESULT resultid="867" eventid="6" status="DSQ" swimtime="00:00:00.00" lane="4" heatid="6001" comment="falscher Start, Gesicht aus dem Wasser (Aufgegeben) nach 130 m">
                  <SPLITS>
                    <SPLIT distance="200" swimtime="00:01:08.25" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="946" eventid="10" status="DSQ" swimtime="00:00:23.12" lane="4" heatid="10002" comment="falscher Start" />
                <RESULT resultid="837" eventid="12" swimtime="00:02:04.66" lane="4" heatid="12005">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:59.73" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="936" eventid="17" swimtime="00:00:24.04" lane="4" heatid="17005" />
                <RESULT resultid="815" eventid="22" swimtime="00:00:52.50" lane="6" heatid="22002" />
                <RESULT resultid="861" eventid="26" swimtime="00:04:23.89" lane="7" heatid="26004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:02.80" />
                    <SPLIT distance="200" swimtime="00:02:13.13" />
                    <SPLIT distance="300" swimtime="00:03:22.35" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="213" birthdate="1978-01-01" gender="M" lastname="Hannemann" firstname="Ronny" license="0">
              <RESULTS>
                <RESULT resultid="803" eventid="2" swimtime="00:00:56.68" lane="6" heatid="2005" />
                <RESULT resultid="888" eventid="8" swimtime="00:00:24.03" lane="8" heatid="8002" />
                <RESULT resultid="937" eventid="17" swimtime="00:00:26.06" lane="2" heatid="17005" />
                <RESULT resultid="813" eventid="22" swimtime="00:01:00.26" lane="8" heatid="22003" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="214" birthdate="2010-01-01" gender="M" lastname="Hochstein" firstname="Jean Paul" license="0">
              <RESULTS>
                <RESULT resultid="804" eventid="2" swimtime="00:01:00.54" lane="6" heatid="2004" />
                <RESULT resultid="948" eventid="10" swimtime="00:00:29.25" lane="2" heatid="10002" />
                <RESULT resultid="840" eventid="12" swimtime="00:02:18.89" lane="5" heatid="12004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:08.74" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="938" eventid="17" swimtime="00:00:26.09" lane="1" heatid="17005" />
                <RESULT resultid="901" eventid="19" swimtime="00:00:28.03" lane="2" heatid="19003" />
                <RESULT resultid="864" eventid="26" swimtime="00:04:52.75" lane="2" heatid="26003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:10.02" />
                    <SPLIT distance="200" swimtime="00:02:25.14" />
                    <SPLIT distance="300" swimtime="00:03:42.11" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="215" birthdate="2010-01-01" gender="M" lastname="Blumenstein" firstname="Einar" license="0">
              <RESULTS>
                <RESULT resultid="806" eventid="2" swimtime="00:01:01.40" lane="7" heatid="2004" />
                <RESULT resultid="842" eventid="12" swimtime="00:02:25.53" lane="6" heatid="12004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:09.31" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="941" eventid="17" swimtime="00:00:28.08" lane="6" heatid="17004" />
                <RESULT resultid="902" eventid="19" swimtime="00:00:27.96" lane="8" heatid="19003" />
                <RESULT resultid="865" eventid="26" swimtime="00:05:35.21" lane="5" heatid="26002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:16.52" />
                    <SPLIT distance="200" swimtime="00:02:46.23" />
                    <SPLIT distance="300" swimtime="00:04:17.35" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="216" birthdate="2009-01-01" gender="F" lastname="Zitzmann" firstname="Annalena" license="0">
              <RESULTS>
                <RESULT resultid="919" eventid="16" swimtime="00:00:22.83" lane="3" heatid="16009" />
                <RESULT resultid="891" eventid="18" swimtime="00:00:27.49" lane="2" heatid="18005" />
                <RESULT resultid="809" eventid="21" swimtime="00:00:52.69" lane="6" heatid="21004" />
                <RESULT resultid="849" eventid="25" swimtime="00:04:41.72" lane="4" heatid="25005">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:03.15" />
                    <SPLIT distance="200" swimtime="00:02:18.11" />
                    <SPLIT distance="300" swimtime="00:03:33.21" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY number="2" gender="F" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="868" eventid="28" swimtime="00:03:29.81" lane="3" heatid="28001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:49.71" />
                    <SPLIT distance="200" swimtime="00:01:44.01" />
                    <SPLIT distance="300" swimtime="00:02:37.46" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="199" number="1" />
                    <RELAYPOSITION athleteid="184" number="2" />
                    <RELAYPOSITION athleteid="216" number="3" />
                    <RELAYPOSITION athleteid="202" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="4" gender="F" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="869" eventid="28" swimtime="00:05:06.86" lane="1" heatid="28001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:20.27" />
                    <SPLIT distance="200" swimtime="00:02:46.37" />
                    <SPLIT distance="300" swimtime="00:03:50.24" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="207" number="1" />
                    <RELAYPOSITION athleteid="192" number="2" />
                    <RELAYPOSITION athleteid="205" number="3" />
                    <RELAYPOSITION athleteid="190" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" gender="F" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="870" eventid="27" swimtime="00:04:47.24" lane="4" heatid="27001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:11.72" />
                    <SPLIT distance="200" swimtime="00:02:20.58" />
                    <SPLIT distance="300" swimtime="00:03:36.22" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="189" number="1" />
                    <RELAYPOSITION athleteid="188" number="2" />
                    <RELAYPOSITION athleteid="206" number="3" />
                    <RELAYPOSITION athleteid="208" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="5" gender="X" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="878" eventid="14" swimtime="00:01:43.08" lane="4" heatid="14001">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="213" number="1" />
                    <RELAYPOSITION athleteid="204" number="2" />
                    <RELAYPOSITION athleteid="185" number="3" />
                    <RELAYPOSITION athleteid="210" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT resultid="871" eventid="29" swimtime="00:03:48.71" lane="6" heatid="29001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:55.89" />
                    <SPLIT distance="200" swimtime="00:01:55.84" />
                    <SPLIT distance="300" swimtime="00:02:58.87" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="213" number="1" />
                    <RELAYPOSITION athleteid="204" number="2" />
                    <RELAYPOSITION athleteid="185" number="3" />
                    <RELAYPOSITION athleteid="210" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="3" gender="M" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="872" eventid="29" swimtime="00:03:59.55" lane="7" heatid="29001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:57.07" />
                    <SPLIT distance="200" swimtime="00:01:55.80" />
                    <SPLIT distance="300" swimtime="00:02:57.16" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="212" number="1" />
                    <RELAYPOSITION athleteid="194" number="2" />
                    <RELAYPOSITION athleteid="214" number="3" />
                    <RELAYPOSITION athleteid="215" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="2" gender="X" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="873" eventid="13" swimtime="00:01:28.93" lane="6" heatid="13003">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="203" number="1" />
                    <RELAYPOSITION athleteid="201" number="2" />
                    <RELAYPOSITION athleteid="211" number="3" />
                    <RELAYPOSITION athleteid="209" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="3" gender="X" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="874" eventid="13" swimtime="00:01:35.53" lane="1" heatid="13003">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="199" number="1" />
                    <RELAYPOSITION athleteid="214" number="2" />
                    <RELAYPOSITION athleteid="202" number="3" />
                    <RELAYPOSITION athleteid="212" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="4" gender="X" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="875" eventid="13" swimtime="00:01:51.58" lane="5" heatid="13002">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="184" number="1" />
                    <RELAYPOSITION athleteid="194" number="2" />
                    <RELAYPOSITION athleteid="215" number="3" />
                    <RELAYPOSITION athleteid="205" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" gender="X" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="876" eventid="13" swimtime="00:02:14.97" lane="4" heatid="13001">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="189" number="1" />
                    <RELAYPOSITION athleteid="188" number="2" />
                    <RELAYPOSITION athleteid="196" number="3" />
                    <RELAYPOSITION athleteid="206" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="6" gender="X" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="877" eventid="13" swimtime="00:02:23.25" lane="5" heatid="13001">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="192" number="1" />
                    <RELAYPOSITION athleteid="191" number="2" />
                    <RELAYPOSITION athleteid="197" number="3" />
                    <RELAYPOSITION athleteid="208" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB name="Tauchsportfreunde Dachau e.V." nation="GER" region="34" code="0">
          <ATHLETES>
            <ATHLETE athleteid="229" birthdate="1969-01-01" gender="M" lastname="Sengpiel" firstname="Alexander" license="0">
              <RESULTS>
                <RESULT resultid="964" eventid="2" swimtime="00:00:59.71" lane="8" heatid="2005" />
                <RESULT resultid="965" eventid="8" swimtime="00:00:23.30" lane="4" heatid="8001" />
                <RESULT resultid="966" eventid="12" swimtime="00:02:14.55" lane="7" heatid="12005">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:04.13" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="967" eventid="20" swimtime="00:11:07.60" lane="3" heatid="20002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:12.43" />
                    <SPLIT distance="200" swimtime="00:02:36.34" />
                    <SPLIT distance="300" swimtime="00:04:02.13" />
                    <SPLIT distance="400" swimtime="00:05:28.93" />
                    <SPLIT distance="500" swimtime="00:06:54.34" />
                    <SPLIT distance="600" swimtime="00:08:22.13" />
                    <SPLIT distance="700" swimtime="00:09:51.62" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="968" eventid="26" swimtime="00:05:15.37" lane="7" heatid="26003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:09.20" />
                    <SPLIT distance="200" swimtime="00:02:35.11" />
                    <SPLIT distance="300" swimtime="00:04:00.45" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="TC Chemie Greiz e.V." nation="GER" region="35" code="0">
          <ATHLETES>
            <ATHLETE athleteid="66" birthdate="2011-01-01" gender="F" lastname="Leonhardt" firstname="Ronja" license="0">
              <RESULTS>
                <RESULT resultid="290" eventid="1" swimtime="00:01:09.38" lane="7" heatid="1005" />
                <RESULT resultid="279" eventid="3" swimtime="00:01:10.47" lane="8" heatid="3004" />
                <RESULT resultid="309" eventid="11" swimtime="00:02:29.69" lane="8" heatid="11006">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:12.78" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="365" eventid="16" swimtime="00:00:31.38" lane="2" heatid="16004" />
                <RESULT resultid="379" eventid="20" swimtime="00:11:07.62" lane="7" heatid="20002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:15.59" />
                    <SPLIT distance="200" swimtime="00:02:41.55" />
                    <SPLIT distance="300" swimtime="00:04:11.54" />
                    <SPLIT distance="400" swimtime="00:05:39.79" />
                    <SPLIT distance="500" swimtime="00:07:03.10" />
                    <SPLIT distance="600" swimtime="00:08:28.97" />
                    <SPLIT distance="700" swimtime="00:09:51.68" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="322" eventid="25" swimtime="00:05:23.05" lane="6" heatid="25004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:14.83" />
                    <SPLIT distance="200" swimtime="00:02:41.21" />
                    <SPLIT distance="300" swimtime="00:04:06.68" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="67" birthdate="2011-01-01" gender="F" lastname="Volger" firstname="Eva" license="0">
              <RESULTS>
                <RESULT resultid="292" eventid="1" swimtime="00:01:12.58" lane="1" heatid="1004" />
                <RESULT resultid="280" eventid="3" swimtime="00:01:14.54" lane="2" heatid="3003" />
                <RESULT resultid="310" eventid="11" swimtime="00:02:45.86" lane="4" heatid="11004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:19.05" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="366" eventid="16" swimtime="00:00:32.81" lane="4" heatid="16003" />
                <RESULT resultid="349" eventid="18" swimtime="00:00:33.42" lane="5" heatid="18003" />
                <RESULT resultid="323" eventid="25" swimtime="00:06:02.88" lane="2" heatid="25003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:23.41" />
                    <SPLIT distance="200" swimtime="00:02:58.61" />
                    <SPLIT distance="300" swimtime="00:04:34.95" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="68" birthdate="2013-01-01" gender="F" lastname="Jutzenka" firstname="Leonie" license="0">
              <RESULTS>
                <RESULT resultid="293" eventid="1" swimtime="00:01:21.86" lane="2" heatid="1003" />
                <RESULT resultid="281" eventid="3" swimtime="00:01:22.76" lane="4" heatid="3002" />
                <RESULT resultid="311" eventid="11" swimtime="00:03:03.12" lane="2" heatid="11003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:26.52" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="367" eventid="16" swimtime="00:00:36.72" lane="7" heatid="16002" />
                <RESULT resultid="350" eventid="18" swimtime="00:00:37.03" lane="1" heatid="18003" />
                <RESULT resultid="356" eventid="23" swimtime="00:00:45.49" lane="1" heatid="23003" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="69" birthdate="2000-01-01" gender="M" lastname="Kupka" firstname="Titus" license="0">
              <RESULTS>
                <RESULT resultid="282" eventid="4" swimtime="00:00:48.92" lane="4" heatid="4003" />
                <RESULT resultid="342" eventid="8" swimtime="00:00:17.01" lane="2" heatid="8004" />
                <RESULT resultid="369" eventid="17" swimtime="00:00:19.59" lane="6" heatid="17008" />
                <RESULT resultid="352" eventid="19" swimtime="00:00:22.09" lane="4" heatid="19004" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="70" birthdate="2008-01-01" gender="M" lastname="Lose" firstname="Fabian" license="0">
              <RESULTS>
                <RESULT resultid="283" eventid="4" swimtime="00:00:58.64" lane="8" heatid="4003" />
                <RESULT resultid="317" eventid="12" swimtime="00:02:12.73" lane="2" heatid="12005">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:03.71" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="353" eventid="19" swimtime="00:00:26.28" lane="6" heatid="19003" />
                <RESULT resultid="326" eventid="26" swimtime="00:04:42.81" lane="4" heatid="26003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:06.37" />
                    <SPLIT distance="200" swimtime="00:02:22.32" />
                    <SPLIT distance="300" swimtime="00:03:35.72" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="71" birthdate="2012-01-01" gender="M" lastname="Sochynskyi" firstname="Vadym" license="0">
              <RESULTS>
                <RESULT resultid="299" eventid="2" swimtime="00:01:16.45" lane="3" heatid="2003" />
                <RESULT resultid="284" eventid="4" swimtime="00:01:09.31" lane="3" heatid="4002" />
                <RESULT resultid="319" eventid="12" swimtime="00:02:34.66" lane="8" heatid="12004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:16.64" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="373" eventid="17" swimtime="00:00:32.42" lane="8" heatid="17004" />
                <RESULT resultid="354" eventid="19" swimtime="00:00:31.03" lane="4" heatid="19002" />
                <RESULT resultid="358" eventid="24" swimtime="00:00:33.03" lane="5" heatid="24002" />
                <RESULT resultid="328" eventid="26" swimtime="00:05:28.26" lane="3" heatid="26002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:16.83" />
                    <SPLIT distance="200" swimtime="00:02:42.69" />
                    <SPLIT distance="300" swimtime="00:04:04.52" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="72" birthdate="2014-01-01" gender="M" lastname="Volger" firstname="Tom" license="0">
              <RESULTS>
                <RESULT resultid="300" eventid="2" swimtime="00:01:17.61" lane="8" heatid="2003" />
                <RESULT resultid="285" eventid="4" swimtime="00:01:20.05" lane="7" heatid="4002" />
                <RESULT resultid="320" eventid="12" swimtime="00:02:48.65" lane="3" heatid="12003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:23.72" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="374" eventid="17" swimtime="00:00:35.38" lane="5" heatid="17002" />
                <RESULT resultid="355" eventid="19" swimtime="00:00:35.66" lane="7" heatid="19002" />
                <RESULT resultid="359" eventid="24" swimtime="00:00:36.49" lane="7" heatid="24002" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="73" birthdate="2005-01-01" gender="F" lastname="Kupka" firstname="Miriam" license="0">
              <RESULTS>
                <RESULT resultid="286" eventid="1" swimtime="00:00:46.00" lane="5" heatid="1012" />
                <RESULT resultid="338" eventid="7" swimtime="00:00:19.65" lane="2" heatid="7005" />
                <RESULT resultid="306" eventid="11" swimtime="00:01:46.41" lane="3" heatid="11010">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:50.56" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="360" eventid="16" swimtime="00:00:20.68" lane="3" heatid="16011" />
                <RESULT resultid="321" eventid="25" swimtime="00:03:50.08" lane="6" heatid="25008">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:53.04" />
                    <SPLIT distance="200" swimtime="00:01:52.04" />
                    <SPLIT distance="300" swimtime="00:02:52.66" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="74" birthdate="2006-01-01" gender="F" lastname="Frauenfelder" firstname="Anneliese" license="0">
              <RESULTS>
                <RESULT resultid="287" eventid="1" swimtime="00:00:48.80" lane="6" heatid="1011" />
                <RESULT resultid="329" eventid="5" swimtime="00:04:16.75" lane="3" heatid="5002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:55.94" />
                    <SPLIT distance="200" swimtime="00:02:01.42" />
                    <SPLIT distance="300" swimtime="00:03:11.53" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="339" eventid="7" swimtime="00:00:21.63" lane="4" heatid="7004" />
                <RESULT resultid="361" eventid="16" swimtime="00:00:22.85" lane="3" heatid="16010" />
                <RESULT resultid="301" eventid="21" swimtime="00:00:47.88" lane="7" heatid="21006" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="75" birthdate="2006-01-01" gender="F" lastname="Löffler" firstname="Johanna" license="0">
              <RESULTS>
                <RESULT resultid="288" eventid="1" swimtime="00:00:52.71" lane="8" heatid="1011" />
                <RESULT resultid="340" eventid="7" swimtime="00:00:21.69" lane="1" heatid="7004" />
                <RESULT resultid="307" eventid="11" swimtime="00:01:59.39" lane="7" heatid="11010">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:58.34" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="362" eventid="16" swimtime="00:00:23.37" lane="6" heatid="16010" />
                <RESULT resultid="346" eventid="18" swimtime="00:00:27.52" lane="6" heatid="18005" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="76" birthdate="2009-01-01" gender="F" lastname="Nauphold" firstname="Celina" license="0">
              <RESULTS>
                <RESULT resultid="289" eventid="1" swimtime="00:00:56.10" lane="2" heatid="1009" />
                <RESULT resultid="341" eventid="7" swimtime="00:00:24.11" lane="3" heatid="7003" />
                <RESULT resultid="363" eventid="16" swimtime="00:00:25.76" lane="8" heatid="16009" />
                <RESULT resultid="347" eventid="18" swimtime="00:00:29.73" lane="3" heatid="18004" />
                <RESULT resultid="303" eventid="21" swimtime="00:00:55.33" lane="5" heatid="21003" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="77" birthdate="2011-01-01" gender="F" lastname="Klar" firstname="Sophia" license="0">
              <RESULTS>
                <RESULT resultid="291" eventid="1" swimtime="00:01:20.49" lane="4" heatid="1004" />
                <RESULT resultid="375" eventid="9" swimtime="00:00:32.40" lane="7" heatid="9002" />
                <RESULT resultid="312" eventid="11" swimtime="00:03:07.66" lane="1" heatid="11003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:31.90" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="364" eventid="16" swimtime="00:00:32.21" lane="1" heatid="16005" />
                <RESULT resultid="380" eventid="20" swimtime="00:13:58.18" lane="1" heatid="20002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:34.09" />
                    <SPLIT distance="200" swimtime="00:03:21.07" />
                    <SPLIT distance="300" swimtime="00:05:10.47" />
                    <SPLIT distance="400" swimtime="00:06:56.83" />
                    <SPLIT distance="500" swimtime="00:08:46.89" />
                    <SPLIT distance="600" swimtime="00:10:38.49" />
                    <SPLIT distance="700" swimtime="00:12:20.99" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="304" eventid="21" swimtime="00:01:21.43" lane="6" heatid="21002" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="78" birthdate="2016-01-01" gender="F" lastname="Volger" firstname="Lea" license="0">
              <RESULTS>
                <RESULT resultid="294" eventid="1" swimtime="00:01:29.55" lane="6" heatid="1002" />
                <RESULT resultid="313" eventid="11" swimtime="00:03:12.83" lane="4" heatid="11001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:37.46" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="368" eventid="16" swimtime="00:00:38.56" lane="1" heatid="16002" />
                <RESULT resultid="351" eventid="18" swimtime="00:00:39.39" lane="8" heatid="18003" />
                <RESULT resultid="357" eventid="23" swimtime="00:00:39.58" lane="7" heatid="23002" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="79" birthdate="2008-01-01" gender="M" lastname="Berger" firstname="Louis" license="0">
              <RESULTS>
                <RESULT resultid="295" eventid="2" swimtime="00:00:44.24" lane="2" heatid="2008" />
                <RESULT resultid="343" eventid="8" status="DSQ" swimtime="00:00:17.61" lane="6" heatid="8003" comment="falscher Start" />
                <RESULT resultid="314" eventid="12" swimtime="00:01:42.21" lane="2" heatid="12007">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:48.22" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="370" eventid="17" swimtime="00:00:19.35" lane="2" heatid="17008" />
                <RESULT resultid="324" eventid="26" swimtime="00:03:47.24" lane="5" heatid="26005">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:50.03" />
                    <SPLIT distance="200" swimtime="00:01:47.15" />
                    <SPLIT distance="300" swimtime="00:02:48.58" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="80" birthdate="1974-01-01" gender="M" lastname="Kühn" firstname="Ronald" license="0">
              <RESULTS>
                <RESULT resultid="296" eventid="2" swimtime="00:00:56.24" lane="6" heatid="2006" />
                <RESULT resultid="344" eventid="8" swimtime="00:00:20.83" lane="6" heatid="8002" />
                <RESULT resultid="316" eventid="12" swimtime="00:02:16.75" lane="5" heatid="12005">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:09.25" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="371" eventid="17" swimtime="00:00:25.46" lane="2" heatid="17006" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="81" birthdate="2009-01-01" gender="M" lastname="Heydel" firstname="Linus" license="0">
              <RESULTS>
                <RESULT resultid="297" eventid="2" swimtime="00:00:52.77" lane="1" heatid="2006" />
                <RESULT resultid="331" eventid="6" swimtime="00:04:37.55" lane="5" heatid="6001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:02.67" />
                    <SPLIT distance="200" swimtime="00:02:15.13" />
                    <SPLIT distance="300" swimtime="00:03:29.85" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="345" eventid="8" swimtime="00:00:21.58" lane="2" heatid="8002" />
                <RESULT resultid="315" eventid="12" swimtime="00:02:03.33" lane="1" heatid="12006">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:58.50" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="372" eventid="17" swimtime="00:00:25.23" lane="3" heatid="17005" />
                <RESULT resultid="377" eventid="20" swimtime="00:09:36.82" lane="7" heatid="20003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:06.11" />
                    <SPLIT distance="200" swimtime="00:02:20.70" />
                    <SPLIT distance="300" swimtime="00:03:36.31" />
                    <SPLIT distance="400" swimtime="00:04:51.26" />
                    <SPLIT distance="500" swimtime="00:06:04.65" />
                    <SPLIT distance="600" swimtime="00:07:19.40" />
                    <SPLIT distance="700" swimtime="00:08:30.38" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="305" eventid="22" swimtime="00:00:55.37" lane="1" heatid="22003" />
                <RESULT resultid="325" eventid="26" swimtime="00:04:29.86" lane="2" heatid="26004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:02.03" />
                    <SPLIT distance="200" swimtime="00:02:13.71" />
                    <SPLIT distance="300" swimtime="00:03:24.58" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="82" birthdate="2011-01-01" gender="M" lastname="Wyczisk" firstname="Johann" license="0">
              <RESULTS>
                <RESULT resultid="298" eventid="2" swimtime="00:01:08.33" lane="1" heatid="2004" />
                <RESULT resultid="376" eventid="10" swimtime="00:00:33.17" lane="7" heatid="10002" />
                <RESULT resultid="318" eventid="12" swimtime="00:02:28.64" lane="2" heatid="12004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:12.01" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="378" eventid="20" swimtime="00:11:57.25" lane="2" heatid="20002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:19.76" />
                    <SPLIT distance="200" swimtime="00:02:51.39" />
                    <SPLIT distance="300" swimtime="00:04:22.04" />
                    <SPLIT distance="400" swimtime="00:05:54.98" />
                    <SPLIT distance="500" swimtime="00:07:28.14" />
                    <SPLIT distance="600" swimtime="00:08:59.48" />
                    <SPLIT distance="700" swimtime="00:10:28.46" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="327" eventid="26" swimtime="00:05:37.69" lane="6" heatid="26003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:12.78" />
                    <SPLIT distance="200" swimtime="00:02:37.74" />
                    <SPLIT distance="300" swimtime="00:04:10.46" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="83" birthdate="2008-01-01" gender="F" lastname="Zschegner" firstname="Lucy" license="0">
              <RESULTS>
                <RESULT resultid="330" eventid="5" status="DNS" swimtime="00:00:00.00" lane="5" heatid="5001" />
                <RESULT resultid="308" eventid="11" status="DNS" swimtime="00:00:00.00" lane="1" heatid="11008" />
                <RESULT resultid="348" eventid="18" status="DNS" swimtime="00:00:00.00" lane="6" heatid="18004" />
                <RESULT resultid="302" eventid="21" status="DNS" swimtime="00:00:00.00" lane="3" heatid="21004" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY number="1" gender="X" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="332" eventid="27" swimtime="00:05:23.48" lane="6" heatid="27001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:17.51" />
                    <SPLIT distance="200" swimtime="00:02:42.66" />
                    <SPLIT distance="300" swimtime="00:04:11.30" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="72" number="1" />
                    <RELAYPOSITION athleteid="68" number="2" />
                    <RELAYPOSITION athleteid="78" number="3" />
                    <RELAYPOSITION athleteid="71" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" gender="F" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="333" eventid="28" swimtime="00:03:29.14" lane="4" heatid="28001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:47.34" />
                    <SPLIT distance="200" swimtime="00:01:44.47" />
                    <SPLIT distance="300" swimtime="00:02:39.52" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="73" number="1" />
                    <RELAYPOSITION athleteid="76" number="2" />
                    <RELAYPOSITION athleteid="75" number="3" />
                    <RELAYPOSITION athleteid="74" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" gender="F" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="334" eventid="28" status="WDR" swimtime="00:00:00.00" lane="7" heatid="28001">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="76" number="1" />
                    <RELAYPOSITION athleteid="67" number="2" />
                    <RELAYPOSITION athleteid="66" number="3" />
                    <RELAYPOSITION athleteid="77" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" gender="X" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="335" eventid="13" swimtime="00:01:21.46" lane="4" heatid="13003">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="73" number="1" />
                    <RELAYPOSITION athleteid="69" number="2" />
                    <RELAYPOSITION athleteid="74" number="3" />
                    <RELAYPOSITION athleteid="79" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" gender="X" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="336" eventid="13" swimtime="00:01:39.87" lane="8" heatid="13003">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="81" number="1" />
                    <RELAYPOSITION athleteid="75" number="2" />
                    <RELAYPOSITION athleteid="70" number="3" />
                    <RELAYPOSITION athleteid="76" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" gender="X" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="337" eventid="13" swimtime="00:02:07.70" lane="6" heatid="13002">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="82" number="1" />
                    <RELAYPOSITION athleteid="71" number="2" />
                    <RELAYPOSITION athleteid="77" number="3" />
                    <RELAYPOSITION athleteid="66" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB name="TC Nautilus Mitterteich e.V." nation="GER" region="34" code="0">
          <ATHLETES>
            <ATHLETE athleteid="227" birthdate="1992-01-01" gender="F" lastname="Schaller" firstname="Christin" license="0">
              <RESULTS>
                <RESULT resultid="958" eventid="1" swimtime="00:01:00.62" lane="6" heatid="1008" />
                <RESULT resultid="959" eventid="11" swimtime="00:02:11.87" lane="5" heatid="11008">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:04.16" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="960" eventid="16" swimtime="00:00:27.46" lane="6" heatid="16006" />
                <RESULT resultid="961" eventid="20" swimtime="00:10:29.65" lane="6" heatid="20003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:11.26" />
                    <SPLIT distance="200" swimtime="00:02:31.43" />
                    <SPLIT distance="300" swimtime="00:03:51.82" />
                    <SPLIT distance="400" swimtime="00:05:12.52" />
                    <SPLIT distance="500" swimtime="00:06:34.24" />
                    <SPLIT distance="600" swimtime="00:07:56.01" />
                    <SPLIT distance="700" swimtime="00:09:15.59" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="962" eventid="21" status="DNS" swimtime="00:00:00.00" lane="7" heatid="21004" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="TC submarin Pößneck" nation="GER" region="35" code="0">
          <ATHLETES>
            <ATHLETE athleteid="234" birthdate="2010-01-01" gender="F" lastname="Matthes" firstname="Sophie" license="0">
              <RESULTS>
                <RESULT resultid="1001" eventid="1" swimtime="00:01:02.09" lane="5" heatid="1007" />
                <RESULT resultid="982" eventid="3" swimtime="00:01:09.44" lane="3" heatid="3004" />
                <RESULT resultid="1096" eventid="9" swimtime="00:00:26.94" lane="5" heatid="9002" />
                <RESULT resultid="1024" eventid="11" swimtime="00:02:26.66" lane="5" heatid="11006">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:10.02" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1083" eventid="16" swimtime="00:00:27.04" lane="1" heatid="16008" />
                <RESULT resultid="1056" eventid="18" swimtime="00:00:29.81" lane="4" heatid="18004" />
                <RESULT resultid="1017" eventid="21" swimtime="00:01:06.14" lane="4" heatid="21002" />
                <RESULT resultid="1037" eventid="25" swimtime="00:05:23.57" lane="4" heatid="25004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:16.48" />
                    <SPLIT distance="200" swimtime="00:02:45.16" />
                    <SPLIT distance="300" swimtime="00:04:11.17" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="235" birthdate="2012-01-01" gender="F" lastname="Kraus" firstname="Letizia Marie" license="0">
              <RESULTS>
                <RESULT resultid="1002" eventid="1" swimtime="00:01:00.92" lane="7" heatid="1007" />
                <RESULT resultid="983" eventid="3" swimtime="00:01:09.05" lane="6" heatid="3004" />
                <RESULT resultid="1023" eventid="11" swimtime="00:02:16.21" lane="3" heatid="11007">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:05.83" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1084" eventid="16" swimtime="00:00:29.04" lane="7" heatid="16007" />
                <RESULT resultid="1055" eventid="18" status="DSQ" swimtime="00:00:31.38" lane="8" heatid="18005" comment="falscher Schwimmstil (keine Arme)" />
                <RESULT resultid="1070" eventid="23" swimtime="00:00:29.71" lane="4" heatid="23004" />
                <RESULT resultid="1036" eventid="25" swimtime="00:04:43.49" lane="7" heatid="25006">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:05.22" />
                    <SPLIT distance="200" swimtime="00:02:19.30" />
                    <SPLIT distance="300" swimtime="00:03:33.28" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="236" birthdate="2011-01-01" gender="F" lastname="Müller" firstname="Emily" license="0">
              <RESULTS>
                <RESULT resultid="1003" eventid="1" swimtime="00:01:08.01" lane="2" heatid="1006" />
                <RESULT resultid="984" eventid="3" swimtime="00:01:11.02" lane="1" heatid="3004" />
                <RESULT resultid="1095" eventid="9" status="DSQ" swimtime="00:00:44.18" lane="5" heatid="9001" comment="Gesich aus dem Wasser (Aufgegeben) nach 8 m" />
                <RESULT resultid="1025" eventid="11" swimtime="00:02:29.24" lane="2" heatid="11005">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:12.40" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1085" eventid="16" swimtime="00:00:30.43" lane="8" heatid="16005" />
                <RESULT resultid="1057" eventid="18" swimtime="00:00:31.83" lane="4" heatid="18003" />
                <RESULT resultid="1013" eventid="21" status="DSQ" swimtime="00:01:21.24" lane="3" heatid="21001" comment="Gesicht aus dem Wasser bei 20m" />
                <RESULT resultid="1038" eventid="25" swimtime="00:05:21.38" lane="4" heatid="25003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:13.82" />
                    <SPLIT distance="200" swimtime="00:02:39.05" />
                    <SPLIT distance="300" swimtime="00:04:05.78" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="237" birthdate="2013-01-01" gender="F" lastname="Huber" firstname="Sina" license="0">
              <RESULTS>
                <RESULT resultid="1004" eventid="1" swimtime="00:01:16.14" lane="5" heatid="1004" />
                <RESULT resultid="985" eventid="3" swimtime="00:01:27.41" lane="7" heatid="3003" />
                <RESULT resultid="1026" eventid="11" swimtime="00:02:45.74" lane="4" heatid="11003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:23.20" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1086" eventid="16" swimtime="00:00:32.38" lane="6" heatid="16004" />
                <RESULT resultid="1059" eventid="18" swimtime="00:00:35.12" lane="6" heatid="18003" />
                <RESULT resultid="1075" eventid="23" swimtime="00:00:37.62" lane="8" heatid="23003" />
                <RESULT resultid="1039" eventid="25" swimtime="00:06:05.31" lane="4" heatid="25002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:27.16" />
                    <SPLIT distance="200" swimtime="00:03:01.69" />
                    <SPLIT distance="300" swimtime="00:04:39.47" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="238" birthdate="2013-01-01" gender="F" lastname="Schmidt" firstname="Ylva" license="0">
              <RESULTS>
                <RESULT resultid="1006" eventid="1" swimtime="00:01:19.18" lane="5" heatid="1003" />
                <RESULT resultid="986" eventid="3" swimtime="00:01:22.72" lane="5" heatid="3002" />
                <RESULT resultid="1028" eventid="11" swimtime="00:02:58.70" lane="6" heatid="11003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:27.93" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1088" eventid="16" swimtime="00:00:34.66" lane="4" heatid="16002" />
                <RESULT resultid="1058" eventid="18" swimtime="00:00:34.15" lane="3" heatid="18003" />
                <RESULT resultid="1071" eventid="23" swimtime="00:00:35.13" lane="5" heatid="23003" />
                <RESULT resultid="1041" eventid="25" swimtime="00:06:05.33" lane="8" heatid="25002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:27.87" />
                    <SPLIT distance="200" swimtime="00:03:02.47" />
                    <SPLIT distance="300" swimtime="00:04:37.85" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="239" birthdate="2013-01-01" gender="F" lastname="Werner" firstname="Zoe" license="0">
              <RESULTS>
                <RESULT resultid="1007" eventid="1" status="DSQ" swimtime="00:01:16.57" lane="3" heatid="1003" comment="falscher Start" />
                <RESULT resultid="987" eventid="3" swimtime="00:01:20.10" lane="3" heatid="3002" />
                <RESULT resultid="1029" eventid="11" swimtime="00:02:48.06" lane="7" heatid="11003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:23.71" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1090" eventid="16" swimtime="00:00:35.22" lane="2" heatid="16002" />
                <RESULT resultid="1062" eventid="18" swimtime="00:00:35.54" lane="5" heatid="18002" />
                <RESULT resultid="1073" eventid="23" swimtime="00:00:38.55" lane="6" heatid="23003" />
                <RESULT resultid="1035" eventid="25" swimtime="00:05:59.00" lane="3" heatid="25001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:26.08" />
                    <SPLIT distance="200" swimtime="00:02:59.89" />
                    <SPLIT distance="300" swimtime="00:04:33.52" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="240" birthdate="2013-01-01" gender="F" lastname="Wolschendorf" firstname="Zoe" license="0">
              <RESULTS>
                <RESULT resultid="1008" eventid="1" swimtime="00:01:20.05" lane="8" heatid="1003" />
                <RESULT resultid="988" eventid="3" swimtime="00:01:23.53" lane="6" heatid="3002" />
                <RESULT resultid="1030" eventid="11" swimtime="00:03:04.38" lane="5" heatid="11002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:25.08" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="241" birthdate="2013-01-01" gender="F" lastname="Dietzel" firstname="Hanna" license="0">
              <RESULTS>
                <RESULT resultid="1009" eventid="1" swimtime="00:01:25.28" lane="5" heatid="1002" />
                <RESULT resultid="989" eventid="3" swimtime="00:01:31.20" lane="2" heatid="3002" />
                <RESULT resultid="1031" eventid="11" swimtime="00:03:19.78" lane="7" heatid="11002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:35.49" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1089" eventid="16" swimtime="00:00:36.04" lane="5" heatid="16002" />
                <RESULT resultid="1061" eventid="18" swimtime="00:00:37.78" lane="4" heatid="18002" />
                <RESULT resultid="1077" eventid="23" swimtime="00:00:46.66" lane="2" heatid="23002" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="242" birthdate="2015-01-01" gender="F" lastname="Knoblich" firstname="Anna" license="0">
              <RESULTS>
                <RESULT resultid="990" eventid="3" swimtime="00:01:51.76" lane="8" heatid="3002" />
                <RESULT resultid="1064" eventid="18" swimtime="00:00:46.61" lane="5" heatid="18001" />
                <RESULT resultid="1078" eventid="23" swimtime="00:00:46.47" lane="4" heatid="23001" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="243" birthdate="2015-01-01" gender="F" lastname="Huber" firstname="Karla" license="0">
              <RESULTS>
                <RESULT resultid="991" eventid="3" swimtime="00:01:32.45" lane="4" heatid="3001" />
                <RESULT resultid="1063" eventid="18" swimtime="00:00:41.72" lane="4" heatid="18001" />
                <RESULT resultid="1072" eventid="23" swimtime="00:00:43.93" lane="3" heatid="23003" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="244" birthdate="2015-01-01" gender="F" lastname="Wolschendorf" firstname="Ella" license="0">
              <RESULTS>
                <RESULT resultid="992" eventid="3" swimtime="00:01:28.02" lane="5" heatid="3001" />
                <RESULT resultid="1021" eventid="11" swimtime="00:03:17.40" lane="2" heatid="11001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:35.08" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="245" birthdate="2014-01-01" gender="F" lastname="Cislak" firstname="Leni" license="0">
              <RESULTS>
                <RESULT resultid="993" eventid="3" swimtime="00:01:41.18" lane="3" heatid="3001" />
                <RESULT resultid="1065" eventid="18" swimtime="00:01:00.65" lane="3" heatid="18001" />
                <RESULT resultid="1074" eventid="23" status="DSQ" swimtime="00:01:20.85" lane="2" heatid="23003" comment="falscher Start" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="246" birthdate="2011-01-01" gender="M" lastname="Rattke" firstname="Carlos" license="0">
              <RESULTS>
                <RESULT resultid="1010" eventid="2" swimtime="00:01:12.60" lane="5" heatid="2003" />
                <RESULT resultid="994" eventid="4" swimtime="00:01:17.59" lane="6" heatid="4002" />
                <RESULT resultid="1097" eventid="10" swimtime="00:00:41.46" lane="3" heatid="10001" />
                <RESULT resultid="1032" eventid="12" swimtime="00:02:44.35" lane="7" heatid="12004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:20.56" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1092" eventid="17" swimtime="00:00:35.80" lane="3" heatid="17003" />
                <RESULT resultid="1066" eventid="19" swimtime="00:00:31.20" lane="5" heatid="19002" />
                <RESULT resultid="1018" eventid="22" swimtime="00:01:28.09" lane="1" heatid="22001" />
                <RESULT resultid="1044" eventid="26" swimtime="00:05:49.16" lane="1" heatid="26003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:24.38" />
                    <SPLIT distance="200" swimtime="00:02:55.01" />
                    <SPLIT distance="300" swimtime="00:04:24.56" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="247" birthdate="2011-01-01" gender="M" lastname="Knoblich" firstname="Paul" license="0">
              <RESULTS>
                <RESULT resultid="1011" eventid="2" swimtime="00:01:10.36" lane="7" heatid="2003" />
                <RESULT resultid="995" eventid="4" swimtime="00:01:19.23" lane="2" heatid="4002" />
                <RESULT resultid="1098" eventid="10" swimtime="00:00:35.10" lane="4" heatid="10001" />
                <RESULT resultid="1033" eventid="12" swimtime="00:02:39.31" lane="4" heatid="12003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:19.96" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1091" eventid="17" status="DSQ" swimtime="00:00:31.73" lane="4" heatid="17003" comment="falscher Start" />
                <RESULT resultid="1099" eventid="20" swimtime="00:12:16.94" lane="3" heatid="20001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:20.43" />
                    <SPLIT distance="200" swimtime="00:02:52.87" />
                    <SPLIT distance="300" swimtime="00:04:27.38" />
                    <SPLIT distance="400" swimtime="00:06:04.37" />
                    <SPLIT distance="500" swimtime="00:07:40.17" />
                    <SPLIT distance="600" swimtime="00:09:17.70" />
                    <SPLIT distance="700" swimtime="00:10:54.89" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1019" eventid="22" swimtime="00:01:26.17" lane="5" heatid="22001" />
                <RESULT resultid="1045" eventid="26" swimtime="00:05:37.34" lane="4" heatid="26002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:22.85" />
                    <SPLIT distance="200" swimtime="00:02:50.03" />
                    <SPLIT distance="300" swimtime="00:04:16.66" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="248" birthdate="2013-01-01" gender="M" lastname="Langlotz" firstname="Lennert" license="0">
              <RESULTS>
                <RESULT resultid="1012" eventid="2" swimtime="00:01:25.81" lane="2" heatid="2002" />
                <RESULT resultid="996" eventid="4" swimtime="00:01:35.38" lane="4" heatid="4001" />
                <RESULT resultid="1034" eventid="12" swimtime="00:03:10.04" lane="4" heatid="12001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:30.59" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="249" birthdate="2016-01-01" gender="M" lastname="Kraus" firstname="Luan" license="0">
              <RESULTS>
                <RESULT resultid="997" eventid="4" swimtime="00:01:36.16" lane="1" heatid="4001" />
                <RESULT resultid="1069" eventid="19" swimtime="00:00:44.79" lane="8" heatid="19002" />
                <RESULT resultid="1080" eventid="24" swimtime="00:00:52.41" lane="5" heatid="24001" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="250" birthdate="2005-01-01" gender="F" lastname="Rattke" firstname="Ninette" license="0">
              <RESULTS>
                <RESULT resultid="998" eventid="1" swimtime="00:00:47.51" lane="2" heatid="1012" />
                <RESULT resultid="1047" eventid="5" swimtime="00:03:59.99" lane="7" heatid="5002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:53.64" />
                    <SPLIT distance="200" swimtime="00:01:55.79" />
                    <SPLIT distance="300" swimtime="00:02:59.83" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1054" eventid="7" swimtime="00:00:20.94" lane="8" heatid="7004" />
                <RESULT resultid="1020" eventid="15" swimtime="00:17:28.85" lane="6" heatid="15002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:59.42" />
                    <SPLIT distance="200" swimtime="00:02:05.77" />
                    <SPLIT distance="300" swimtime="00:03:15.57" />
                    <SPLIT distance="400" swimtime="00:04:25.51" />
                    <SPLIT distance="500" swimtime="00:05:36.52" />
                    <SPLIT distance="600" swimtime="00:06:47.36" />
                    <SPLIT distance="700" swimtime="00:07:58.98" />
                    <SPLIT distance="800" swimtime="00:09:09.88" />
                    <SPLIT distance="900" swimtime="00:10:21.53" />
                    <SPLIT distance="1000" swimtime="00:11:33.22" />
                    <SPLIT distance="1100" swimtime="00:12:45.73" />
                    <SPLIT distance="1200" swimtime="00:13:57.53" />
                    <SPLIT distance="1300" swimtime="00:15:09.90" />
                    <SPLIT distance="1400" swimtime="00:16:22.85" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1100" eventid="20" swimtime="00:08:48.84" lane="1" heatid="20004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:55.65" />
                    <SPLIT distance="200" swimtime="00:02:02.00" />
                    <SPLIT distance="300" swimtime="00:03:10.00" />
                    <SPLIT distance="400" swimtime="00:04:20.68" />
                    <SPLIT distance="500" swimtime="00:05:30.95" />
                    <SPLIT distance="600" swimtime="00:06:40.16" />
                    <SPLIT distance="700" swimtime="00:07:47.45" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1015" eventid="21" swimtime="00:00:46.41" lane="1" heatid="21006" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="251" birthdate="2007-01-01" gender="F" lastname="Näther" firstname="Emilia" license="0">
              <RESULTS>
                <RESULT resultid="999" eventid="1" swimtime="00:00:50.06" lane="7" heatid="1011" />
                <RESULT resultid="1048" eventid="5" swimtime="00:04:00.18" lane="8" heatid="5002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:53.32" />
                    <SPLIT distance="200" swimtime="00:01:54.91" />
                    <SPLIT distance="300" swimtime="00:03:00.50" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1053" eventid="7" swimtime="00:00:19.61" lane="1" heatid="7005" />
                <RESULT resultid="1022" eventid="11" swimtime="00:01:49.48" lane="2" heatid="11010">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:51.88" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1082" eventid="16" swimtime="00:00:20.50" lane="5" heatid="16011" />
                <RESULT resultid="1016" eventid="21" swimtime="00:00:46.85" lane="5" heatid="21005" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="252" birthdate="2005-01-01" gender="F" lastname="Heinze" firstname="Charlotte" license="0">
              <RESULTS>
                <RESULT resultid="1000" eventid="1" swimtime="00:00:49.44" lane="1" heatid="1011" />
                <RESULT resultid="1046" eventid="5" swimtime="00:03:58.54" lane="2" heatid="5002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:56.60" />
                    <SPLIT distance="200" swimtime="00:01:57.92" />
                    <SPLIT distance="300" swimtime="00:03:00.43" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1052" eventid="7" swimtime="00:00:18.98" lane="6" heatid="7005" />
                <RESULT resultid="1014" eventid="21" swimtime="00:00:43.51" lane="6" heatid="21006" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="253" birthdate="2013-01-01" gender="F" lastname="Trunk" firstname="Mila" license="0">
              <RESULTS>
                <RESULT resultid="1005" eventid="1" swimtime="00:01:20.41" lane="8" heatid="1004" />
                <RESULT resultid="1027" eventid="11" swimtime="00:02:59.64" lane="3" heatid="11003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:26.65" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1087" eventid="16" swimtime="00:00:33.96" lane="8" heatid="16003" />
                <RESULT resultid="1060" eventid="18" swimtime="00:00:35.94" lane="7" heatid="18003" />
                <RESULT resultid="1076" eventid="23" swimtime="00:00:38.51" lane="3" heatid="23002" />
                <RESULT resultid="1040" eventid="25" swimtime="00:06:00.76" lane="7" heatid="25002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:26.35" />
                    <SPLIT distance="200" swimtime="00:03:00.11" />
                    <SPLIT distance="300" swimtime="00:04:27.63" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="254" birthdate="2013-01-01" gender="M" lastname="Dommler" firstname="Fabrice" license="0">
              <RESULTS>
                <RESULT resultid="1093" eventid="17" swimtime="00:00:36.50" lane="7" heatid="17003" />
                <RESULT resultid="1067" eventid="19" swimtime="00:00:39.28" lane="2" heatid="19002" />
                <RESULT resultid="1079" eventid="24" status="DSQ" swimtime="00:00:44.37" lane="1" heatid="24002" comment="falscher Schwimmstil (Beinwechselschlag) bei 25m" />
                <RESULT resultid="1042" eventid="26" swimtime="00:06:21.51" lane="6" heatid="26001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:26.65" />
                    <SPLIT distance="200" swimtime="00:03:05.25" />
                    <SPLIT distance="300" swimtime="00:04:38.17" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="255" birthdate="2013-01-01" gender="M" lastname="Röser" firstname="Toni" license="0">
              <RESULTS>
                <RESULT resultid="1094" eventid="17" swimtime="00:00:36.10" lane="2" heatid="17002" />
                <RESULT resultid="1068" eventid="19" swimtime="00:00:40.40" lane="1" heatid="19002" />
                <RESULT resultid="1081" eventid="24" swimtime="00:00:51.85" lane="7" heatid="24001" />
                <RESULT resultid="1043" eventid="26" swimtime="00:06:21.65" lane="7" heatid="26001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:29.83" />
                    <SPLIT distance="200" swimtime="00:03:09.13" />
                    <SPLIT distance="300" swimtime="00:04:50.58" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY number="1" gender="X" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="1049" eventid="27" swimtime="00:05:07.93" lane="5" heatid="27001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:20.25" />
                    <SPLIT distance="200" swimtime="00:02:37.04" />
                    <SPLIT distance="300" swimtime="00:04:02.61" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="253" number="1" />
                    <RELAYPOSITION athleteid="237" number="2" />
                    <RELAYPOSITION athleteid="254" number="3" />
                    <RELAYPOSITION athleteid="235" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" gender="X" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="1050" eventid="13" swimtime="00:02:01.52" lane="3" heatid="13002">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="236" number="1" />
                    <RELAYPOSITION athleteid="246" number="2" />
                    <RELAYPOSITION athleteid="247" number="3" />
                    <RELAYPOSITION athleteid="234" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" gender="X" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="1051" eventid="13" swimtime="00:02:14.03" lane="1" heatid="13002">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="239" number="1" />
                    <RELAYPOSITION athleteid="237" number="2" />
                    <RELAYPOSITION athleteid="253" number="3" />
                    <RELAYPOSITION athleteid="235" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" gender="X" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="1101" eventid="13" swimtime="00:02:34.05" lane="8" heatid="13002">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="241" number="1" />
                    <RELAYPOSITION athleteid="243" number="2" />
                    <RELAYPOSITION athleteid="248" number="3" />
                    <RELAYPOSITION athleteid="238" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" gender="X" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="1103" eventid="27" swimtime="00:05:31.43" lane="3" heatid="27001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:25.19" />
                    <SPLIT distance="200" swimtime="00:02:45.32" />
                    <SPLIT distance="300" swimtime="00:04:11.26" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="255" number="1" />
                    <RELAYPOSITION athleteid="239" number="2" />
                    <RELAYPOSITION athleteid="241" number="3" />
                    <RELAYPOSITION athleteid="238" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" gender="X" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="1104" eventid="27" swimtime="00:07:35.81" lane="7" heatid="27001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:02:22.89" />
                    <SPLIT distance="200" swimtime="00:04:17.19" />
                    <SPLIT distance="300" swimtime="00:05:51.90" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="245" number="1" />
                    <RELAYPOSITION athleteid="242" number="2" />
                    <RELAYPOSITION athleteid="249" number="3" />
                    <RELAYPOSITION athleteid="243" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB name="TSC Schwandorf e.V." nation="GER" region="34" code="0">
          <ATHLETES>
            <ATHLETE athleteid="30" birthdate="2004-01-01" gender="F" lastname="Kohler" firstname="Nina" license="0">
              <RESULTS>
                <RESULT resultid="122" eventid="1" swimtime="00:00:43.69" lane="4" heatid="1012" />
                <RESULT resultid="138" eventid="7" swimtime="00:00:17.90" lane="4" heatid="7005" />
                <RESULT resultid="132" eventid="11" swimtime="00:01:37.63" lane="4" heatid="11010">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:46.87" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="141" eventid="16" status="DSQ" swimtime="00:00:19.67" lane="4" heatid="16011" comment="15m nach Start übertaucht" />
                <RESULT resultid="127" eventid="21" swimtime="00:00:41.08" lane="4" heatid="21006" />
                <RESULT resultid="137" eventid="25" swimtime="00:03:41.40" lane="7" heatid="25008">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:52.63" />
                    <SPLIT distance="200" swimtime="00:01:49.74" />
                    <SPLIT distance="300" swimtime="00:02:47.54" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="32" birthdate="2010-01-01" gender="F" lastname="Seitz" firstname="Melina" license="0">
              <RESULTS>
                <RESULT resultid="124" eventid="1" swimtime="00:00:58.50" lane="8" heatid="1008" />
                <RESULT resultid="134" eventid="11" swimtime="00:02:16.73" lane="6" heatid="11004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:04.80" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="142" eventid="16" swimtime="00:00:25.71" lane="6" heatid="16007" />
                <RESULT resultid="128" eventid="21" swimtime="00:01:00.20" lane="1" heatid="21003" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="33" birthdate="2011-01-01" gender="F" lastname="Maget" firstname="Matilda" license="0">
              <RESULTS>
                <RESULT resultid="125" eventid="1" swimtime="00:01:05.20" lane="7" heatid="1006" />
                <RESULT resultid="133" eventid="11" swimtime="00:02:27.38" lane="2" heatid="11004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:10.07" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="143" eventid="16" swimtime="00:00:28.24" lane="4" heatid="16005" />
                <RESULT resultid="129" eventid="21" swimtime="00:01:16.68" lane="3" heatid="21002" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="34" birthdate="2007-01-01" gender="F" lastname="Böhner" firstname="Madeleine" license="0">
              <RESULTS>
                <RESULT resultid="126" eventid="1" swimtime="00:01:08.92" lane="3" heatid="1005" />
                <RESULT resultid="135" eventid="11" swimtime="00:02:35.22" lane="7" heatid="11004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:11.92" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="144" eventid="16" swimtime="00:00:30.62" lane="5" heatid="16004" />
                <RESULT resultid="130" eventid="21" status="DSQ" swimtime="00:01:13.13" lane="2" heatid="21002" comment="falscher Start" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="35" birthdate="2007-01-01" gender="F" lastname="Rödl" firstname="Emily" license="0">
              <RESULTS>
                <RESULT resultid="146" eventid="1" swimtime="00:00:47.75" lane="8" heatid="1012" />
                <RESULT resultid="139" eventid="7" swimtime="00:00:19.98" lane="6" heatid="7004" />
                <RESULT resultid="131" eventid="15" swimtime="00:16:00.01" lane="3" heatid="15002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:57.81" />
                    <SPLIT distance="200" swimtime="00:02:02.36" />
                    <SPLIT distance="300" swimtime="00:03:07.82" />
                    <SPLIT distance="400" swimtime="00:04:14.24" />
                    <SPLIT distance="500" swimtime="00:05:20.15" />
                    <SPLIT distance="600" swimtime="00:06:26.39" />
                    <SPLIT distance="700" swimtime="00:07:32.18" />
                    <SPLIT distance="800" swimtime="00:08:36.81" />
                    <SPLIT distance="900" swimtime="00:09:41.50" />
                    <SPLIT distance="1000" swimtime="00:10:46.04" />
                    <SPLIT distance="1100" swimtime="00:11:49.89" />
                    <SPLIT distance="1200" swimtime="00:12:54.62" />
                    <SPLIT distance="1300" swimtime="00:13:59.42" />
                    <SPLIT distance="1400" swimtime="00:15:02.23" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="140" eventid="18" swimtime="00:00:25.29" lane="3" heatid="18005" />
                <RESULT resultid="145" eventid="20" swimtime="00:08:18.30" lane="6" heatid="20004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:57.43" />
                    <SPLIT distance="200" swimtime="00:02:01.04" />
                    <SPLIT distance="300" swimtime="00:03:05.47" />
                    <SPLIT distance="400" swimtime="00:04:09.65" />
                    <SPLIT distance="500" swimtime="00:05:13.79" />
                    <SPLIT distance="600" swimtime="00:06:18.41" />
                    <SPLIT distance="700" swimtime="00:07:21.06" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="136" eventid="25" swimtime="00:03:59.72" lane="2" heatid="25008">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:56.98" />
                    <SPLIT distance="200" swimtime="00:02:00.55" />
                    <SPLIT distance="300" swimtime="00:03:02.71" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="TSC Weimar e.V." nation="GER" region="35" code="0">
          <ATHLETES>
            <ATHLETE athleteid="98" birthdate="2014-01-01" gender="F" lastname="Rudolph" firstname="Amelie" license="0">
              <RESULTS>
                <RESULT resultid="423" eventid="1" swimtime="00:01:41.30" lane="3" heatid="1001" />
                <RESULT resultid="416" eventid="3" swimtime="00:01:40.12" lane="6" heatid="3001" />
                <RESULT resultid="463" eventid="11" swimtime="00:03:16.68" lane="3" heatid="11001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:35.34" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="525" eventid="16" swimtime="00:00:38.88" lane="6" heatid="16001" />
                <RESULT resultid="499" eventid="18" swimtime="00:00:44.48" lane="2" heatid="18002" />
                <RESULT resultid="510" eventid="23" swimtime="00:00:43.11" lane="5" heatid="23001" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="99" birthdate="2010-01-01" gender="F" lastname="Pontes" firstname="Lena" license="0">
              <RESULTS>
                <RESULT resultid="427" eventid="1" swimtime="00:01:03.10" lane="1" heatid="1007" />
                <RESULT resultid="417" eventid="3" swimtime="00:01:08.19" lane="6" heatid="3003" />
                <RESULT resultid="459" eventid="11" swimtime="00:02:34.66" lane="5" heatid="11005">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:16.17" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="518" eventid="16" swimtime="00:00:27.26" lane="5" heatid="16007" />
                <RESULT resultid="497" eventid="18" swimtime="00:00:29.61" lane="7" heatid="18004" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="100" birthdate="2011-01-01" gender="F" lastname="Hüttig" firstname="Maline" license="0">
              <RESULTS>
                <RESULT resultid="429" eventid="1" swimtime="00:01:08.53" lane="8" heatid="1006" />
                <RESULT resultid="418" eventid="3" swimtime="00:01:18.52" lane="8" heatid="3003" />
                <RESULT resultid="460" eventid="11" swimtime="00:02:56.18" lane="8" heatid="11004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:23.38" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="519" eventid="16" swimtime="00:00:28.43" lane="3" heatid="16006" />
                <RESULT resultid="498" eventid="18" swimtime="00:00:32.71" lane="1" heatid="18004" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="101" birthdate="2007-01-01" gender="M" lastname="Röthlich" firstname="Finn" license="0">
              <RESULTS>
                <RESULT resultid="419" eventid="4" swimtime="00:00:54.07" lane="6" heatid="4003" />
                <RESULT resultid="492" eventid="8" status="DSQ" swimtime="00:00:20.34" lane="1" heatid="8003" comment="falscher Start" />
                <RESULT resultid="963" eventid="19" swimtime="00:00:23.72" lane="2" heatid="19004" />
                <RESULT resultid="451" eventid="22" swimtime="00:00:50.14" lane="2" heatid="22003" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="102" birthdate="2006-01-01" gender="M" lastname="Hauser" firstname="Theo" license="0">
              <RESULTS>
                <RESULT resultid="435" eventid="2" swimtime="00:00:44.48" lane="3" heatid="2007" />
                <RESULT resultid="420" eventid="4" swimtime="00:00:50.69" lane="2" heatid="4003" />
                <RESULT resultid="490" eventid="8" swimtime="00:00:18.47" lane="2" heatid="8003" />
                <RESULT resultid="527" eventid="17" swimtime="00:00:19.68" lane="5" heatid="17007" />
                <RESULT resultid="500" eventid="19" swimtime="00:00:22.44" lane="6" heatid="19004" />
                <RESULT resultid="450" eventid="22" swimtime="00:00:45.74" lane="6" heatid="22003" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="103" birthdate="1968-01-01" gender="M" lastname="Klabunde" firstname="Sven" license="0">
              <RESULTS>
                <RESULT resultid="421" eventid="4" swimtime="00:00:57.30" lane="1" heatid="4003" />
                <RESULT resultid="493" eventid="8" swimtime="00:00:21.90" lane="3" heatid="8001" />
                <RESULT resultid="505" eventid="19" swimtime="00:00:26.11" lane="3" heatid="19003" />
                <RESULT resultid="452" eventid="22" swimtime="00:00:49.34" lane="7" heatid="22002" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="104" birthdate="1956-01-01" gender="M" lastname="Scheffzük" firstname="Olaf" license="0">
              <RESULTS>
                <RESULT resultid="440" eventid="2" swimtime="00:01:01.19" lane="3" heatid="2004" />
                <RESULT resultid="422" eventid="4" swimtime="00:01:06.29" lane="5" heatid="4002" />
                <RESULT resultid="494" eventid="8" swimtime="00:00:30.52" lane="1" heatid="8001" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="105" birthdate="2002-01-01" gender="F" lastname="Kluge" firstname="Paula" license="0">
              <RESULTS>
                <RESULT resultid="424" eventid="1" swimtime="00:00:49.84" lane="3" heatid="1011" />
                <RESULT resultid="472" eventid="5" swimtime="00:04:53.22" lane="1" heatid="5002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:03.53" />
                    <SPLIT distance="200" swimtime="00:02:23.37" />
                    <SPLIT distance="300" swimtime="00:03:41.39" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="483" eventid="7" swimtime="00:00:21.83" lane="3" heatid="7005" />
                <RESULT resultid="516" eventid="16" status="DNS" swimtime="00:00:00.00" lane="1" heatid="16011" />
                <RESULT resultid="444" eventid="21" status="DNS" swimtime="00:00:00.00" lane="3" heatid="21006" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="106" birthdate="2002-01-01" gender="F" lastname="Klabunde" firstname="Lotte" license="0">
              <RESULTS>
                <RESULT resultid="425" eventid="1" swimtime="00:00:48.29" lane="2" heatid="1011" />
                <RESULT resultid="485" eventid="7" swimtime="00:00:19.43" lane="7" heatid="7004" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="107" birthdate="1971-01-01" gender="F" lastname="Klabunde" firstname="Monique" license="0">
              <RESULTS>
                <RESULT resultid="426" eventid="1" swimtime="00:00:53.74" lane="5" heatid="1009" />
                <RESULT resultid="486" eventid="7" swimtime="00:00:23.36" lane="1" heatid="7002" />
                <RESULT resultid="457" eventid="11" swimtime="00:02:01.61" lane="8" heatid="11009">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:58.38" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="469" eventid="25" swimtime="00:04:17.18" lane="8" heatid="25007">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:00.06" />
                    <SPLIT distance="200" swimtime="00:02:06.21" />
                    <SPLIT distance="300" swimtime="00:03:12.65" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="108" birthdate="2010-01-01" gender="F" lastname="Seyfarth" firstname="Annie" license="0">
              <RESULTS>
                <RESULT resultid="428" eventid="1" swimtime="00:01:07.02" lane="4" heatid="1006" />
                <RESULT resultid="458" eventid="11" swimtime="00:02:12.84" lane="3" heatid="11006">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:04.83" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="520" eventid="16" swimtime="00:00:29.06" lane="2" heatid="16006" />
                <RESULT resultid="538" eventid="20" swimtime="00:11:19.26" lane="5" heatid="20001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:12.36" />
                    <SPLIT distance="200" swimtime="00:02:41.12" />
                    <SPLIT distance="300" swimtime="00:04:10.19" />
                    <SPLIT distance="400" swimtime="00:05:40.31" />
                    <SPLIT distance="500" swimtime="00:07:08.67" />
                    <SPLIT distance="600" swimtime="00:08:37.15" />
                    <SPLIT distance="700" swimtime="00:09:58.87" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="470" eventid="25" swimtime="00:05:06.99" lane="3" heatid="25004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:09.74" />
                    <SPLIT distance="200" swimtime="00:02:34.36" />
                    <SPLIT distance="300" swimtime="00:03:57.27" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="109" birthdate="2012-01-01" gender="F" lastname="Linne" firstname="Nora" license="0">
              <RESULTS>
                <RESULT resultid="430" eventid="1" swimtime="00:01:27.88" lane="3" heatid="1002" />
                <RESULT resultid="462" eventid="11" status="DSQ" swimtime="00:03:03.80" lane="2" heatid="11002" comment="falscher Start">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:30.06" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="523" eventid="16" status="DNS" swimtime="00:00:00.00" lane="8" heatid="16002" />
                <RESULT resultid="513" eventid="23" status="DNS" swimtime="00:00:00.00" lane="7" heatid="23003" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="110" birthdate="2013-01-01" gender="F" lastname="Erfurt" firstname="Marit" license="0">
              <RESULTS>
                <RESULT resultid="431" eventid="1" swimtime="00:01:23.63" lane="2" heatid="1002" />
                <RESULT resultid="461" eventid="11" swimtime="00:03:12.49" lane="6" heatid="11002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:32.46" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="524" eventid="16" swimtime="00:00:39.27" lane="4" heatid="16001" />
                <RESULT resultid="512" eventid="23" status="DSQ" swimtime="00:00:44.13" lane="4" heatid="23003" comment="falscher Start" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="111" birthdate="2012-01-01" gender="F" lastname="Gollhardt" firstname="Fridoline" license="0">
              <RESULTS>
                <RESULT resultid="432" eventid="1" swimtime="00:01:14.84" lane="5" heatid="1001" />
                <RESULT resultid="456" eventid="11" swimtime="00:02:49.88" lane="6" heatid="11001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:22.83" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="521" eventid="16" status="DSQ" swimtime="00:00:32.83" lane="3" heatid="16003" comment="falscher Start" />
                <RESULT resultid="511" eventid="23" swimtime="00:00:35.71" lane="1" heatid="23004" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="112" birthdate="2005-01-01" gender="M" lastname="Linne" firstname="Georg" license="0">
              <RESULTS>
                <RESULT resultid="433" eventid="2" swimtime="00:00:43.57" lane="7" heatid="2008" />
                <RESULT resultid="475" eventid="6" swimtime="00:03:12.38" lane="5" heatid="6002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:44.26" />
                    <SPLIT distance="200" swimtime="00:01:32.63" />
                    <SPLIT distance="300" swimtime="00:02:22.39" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="487" eventid="8" swimtime="00:00:17.42" lane="8" heatid="8004" />
                <RESULT resultid="464" eventid="12" swimtime="00:01:38.34" lane="6" heatid="12007">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:46.71" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="504" eventid="19" swimtime="00:00:23.60" lane="8" heatid="19004" />
                <RESULT resultid="446" eventid="22" swimtime="00:00:38.80" lane="5" heatid="22004" />
                <RESULT resultid="471" eventid="26" swimtime="00:03:34.08" lane="3" heatid="26005">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:46.94" />
                    <SPLIT distance="200" swimtime="00:01:40.73" />
                    <SPLIT distance="300" swimtime="00:02:37.38" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="113" birthdate="2004-01-01" gender="M" lastname="Haufe" firstname="Elias" license="0">
              <RESULTS>
                <RESULT resultid="434" eventid="2" swimtime="00:00:44.38" lane="8" heatid="2008" />
                <RESULT resultid="488" eventid="8" swimtime="00:00:15.97" lane="4" heatid="8003" />
                <RESULT resultid="526" eventid="17" swimtime="00:00:18.71" lane="7" heatid="17008" />
                <RESULT resultid="502" eventid="19" swimtime="00:00:22.77" lane="1" heatid="19004" />
                <RESULT resultid="448" eventid="22" swimtime="00:00:43.73" lane="5" heatid="22003" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="114" birthdate="2004-01-01" gender="M" lastname="Röthlich" firstname="Nils" license="0">
              <RESULTS>
                <RESULT resultid="436" eventid="2" swimtime="00:00:47.03" lane="6" heatid="2007" />
                <RESULT resultid="491" eventid="8" swimtime="00:00:18.96" lane="7" heatid="8003" />
                <RESULT resultid="529" eventid="17" swimtime="00:00:20.79" lane="2" heatid="17007" />
                <RESULT resultid="501" eventid="19" swimtime="00:00:24.42" lane="7" heatid="19004" />
                <RESULT resultid="449" eventid="22" swimtime="00:00:45.14" lane="3" heatid="22003" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="115" birthdate="2008-01-01" gender="M" lastname="Kraft" firstname="Simon" license="0">
              <RESULTS>
                <RESULT resultid="437" eventid="2" status="DNS" swimtime="00:00:00.00" lane="2" heatid="2007" />
                <RESULT resultid="528" eventid="17" status="DNS" swimtime="00:00:00.00" lane="6" heatid="17007" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="116" birthdate="2011-01-01" gender="M" lastname="Bellmann" firstname="Lennart" license="0">
              <RESULTS>
                <RESULT resultid="438" eventid="2" swimtime="00:00:57.43" lane="1" heatid="2005" />
                <RESULT resultid="537" eventid="10" swimtime="00:00:28.69" lane="6" heatid="10002" />
                <RESULT resultid="466" eventid="12" swimtime="00:02:12.16" lane="3" heatid="12004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:07.48" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="531" eventid="17" swimtime="00:00:24.58" lane="6" heatid="17005" />
                <RESULT resultid="454" eventid="22" swimtime="00:01:00.24" lane="3" heatid="22001" />
                <RESULT resultid="976" eventid="26" swimtime="00:04:35.04" lane="3" heatid="26003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:07.01" />
                    <SPLIT distance="200" swimtime="00:02:20.02" />
                    <SPLIT distance="300" swimtime="00:03:30.20" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="117" birthdate="2010-01-01" gender="M" lastname="Bellmann" firstname="Arvid" license="0">
              <RESULTS>
                <RESULT resultid="439" eventid="2" swimtime="00:00:59.02" lane="4" heatid="2004" />
                <RESULT resultid="474" eventid="6" swimtime="00:05:19.40" lane="3" heatid="6001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:12.35" />
                    <SPLIT distance="200" swimtime="00:02:32.29" />
                    <SPLIT distance="300" swimtime="00:04:05.17" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="536" eventid="10" swimtime="00:00:25.76" lane="3" heatid="10002" />
                <RESULT resultid="532" eventid="17" status="DSQ" swimtime="00:00:30.48" lane="7" heatid="17005" comment="Tauchzüge (45-46m)" />
                <RESULT resultid="506" eventid="19" swimtime="00:00:29.35" lane="7" heatid="19003" />
                <RESULT resultid="453" eventid="22" swimtime="00:00:59.08" lane="1" heatid="22002" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="118" birthdate="2009-01-01" gender="M" lastname="Klabunde" firstname="Kalle" license="0">
              <RESULTS>
                <RESULT resultid="441" eventid="2" swimtime="00:01:03.20" lane="2" heatid="2004" />
                <RESULT resultid="465" eventid="12" swimtime="00:02:28.51" lane="4" heatid="12004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:10.45" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="533" eventid="17" swimtime="00:00:27.99" lane="3" heatid="17004" />
                <RESULT resultid="508" eventid="19" swimtime="00:00:32.29" lane="6" heatid="19002" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="119" birthdate="1960-01-01" gender="M" lastname="Kaleta" firstname="Bernd" license="0">
              <RESULTS>
                <RESULT resultid="442" eventid="2" swimtime="00:01:12.75" lane="4" heatid="2003" />
                <RESULT resultid="495" eventid="8" swimtime="00:00:33.15" lane="8" heatid="8001" />
                <RESULT resultid="534" eventid="17" swimtime="00:00:31.31" lane="1" heatid="17004" />
                <RESULT resultid="455" eventid="22" swimtime="00:01:21.16" lane="2" heatid="22001" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="120" birthdate="2014-01-01" gender="M" lastname="Schmeißer" firstname="Edwin" license="0">
              <RESULTS>
                <RESULT resultid="443" eventid="2" swimtime="00:01:31.08" lane="4" heatid="2001" />
                <RESULT resultid="467" eventid="12" swimtime="00:03:20.96" lane="3" heatid="12002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:39.95" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="535" eventid="17" swimtime="00:00:44.06" lane="4" heatid="17001" />
                <RESULT resultid="509" eventid="19" swimtime="00:00:42.84" lane="6" heatid="19001" />
                <RESULT resultid="515" eventid="24" swimtime="00:00:48.84" lane="6" heatid="24001" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="128" birthdate="2012-01-01" gender="F" lastname="Riemann" firstname="Ada" license="0">
              <RESULTS>
                <RESULT resultid="522" eventid="16" swimtime="00:00:37.96" lane="6" heatid="16002" />
                <RESULT resultid="514" eventid="23" swimtime="00:00:44.16" lane="5" heatid="23002" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="228" birthdate="1967-01-01" gender="M" lastname="Wurzbacher" firstname="Markus" license="0" />
          </ATHLETES>
          <RELAYS>
            <RELAY number="1" gender="M" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="477" eventid="29" swimtime="00:03:03.95" lane="5" heatid="29001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:43.25" />
                    <SPLIT distance="200" swimtime="00:01:35.57" />
                    <SPLIT distance="300" swimtime="00:02:20.99" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="112" number="1" />
                    <RELAYPOSITION athleteid="101" number="2" />
                    <RELAYPOSITION athleteid="114" number="3" />
                    <RELAYPOSITION athleteid="113" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" gender="X" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="479" eventid="29" swimtime="00:04:08.97" lane="2" heatid="29001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:53.87" />
                    <SPLIT distance="200" swimtime="00:01:54.81" />
                    <SPLIT distance="300" swimtime="00:03:08.94" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="107" number="1" />
                    <RELAYPOSITION athleteid="228" number="2" />
                    <RELAYPOSITION athleteid="119" number="3" />
                    <RELAYPOSITION athleteid="103" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" gender="X" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="480" eventid="13" swimtime="00:01:24.36" lane="2" heatid="13003">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="113" number="1" />
                    <RELAYPOSITION athleteid="106" number="2" />
                    <RELAYPOSITION athleteid="114" number="3" />
                    <RELAYPOSITION athleteid="105" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" gender="X" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="481" eventid="13" swimtime="00:01:47.55" lane="4" heatid="13002">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="117" number="1" />
                    <RELAYPOSITION athleteid="100" number="2" />
                    <RELAYPOSITION athleteid="99" number="3" />
                    <RELAYPOSITION athleteid="116" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" gender="X" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="482" eventid="14" swimtime="00:01:49.01" lane="5" heatid="14001">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="107" number="1" />
                    <RELAYPOSITION athleteid="104" number="2" />
                    <RELAYPOSITION athleteid="119" number="3" />
                    <RELAYPOSITION athleteid="103" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB name="TSG Schwäbisch Hall" nation="GER" region="32" code="0">
          <ATHLETES>
            <ATHLETE athleteid="29" birthdate="1967-01-01" gender="M" lastname="Lochstampfer" firstname="Gunter" license="0">
              <RESULTS>
                <RESULT resultid="118" eventid="2" swimtime="00:00:56.57" lane="2" heatid="2005" />
                <RESULT resultid="117" eventid="4" swimtime="00:00:55.75" lane="7" heatid="4003" />
                <RESULT resultid="119" eventid="8" swimtime="00:00:24.20" lane="5" heatid="8001" />
                <RESULT resultid="121" eventid="17" swimtime="00:00:25.19" lane="5" heatid="17005" />
                <RESULT resultid="120" eventid="19" swimtime="00:00:25.03" lane="4" heatid="19003" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="TSG TU Ilmenau 56 e.V." nation="GER" region="35" code="0">
          <ATHLETES>
            <ATHLETE athleteid="170" birthdate="1999-01-01" gender="F" lastname="Fischer" firstname="Ernestine" license="0">
              <RESULTS>
                <RESULT resultid="697" eventid="1" swimtime="00:00:53.63" lane="1" heatid="1012" />
                <RESULT resultid="977" eventid="5" swimtime="00:04:15.77" lane="6" heatid="5002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:55.29" />
                    <SPLIT distance="200" swimtime="00:02:01.64" />
                    <SPLIT distance="300" swimtime="00:03:12.01" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="741" eventid="7" swimtime="00:00:19.48" lane="5" heatid="7005" />
                <RESULT resultid="748" eventid="16" swimtime="00:00:21.67" lane="2" heatid="16011" />
                <RESULT resultid="710" eventid="21" swimtime="00:00:45.06" lane="5" heatid="21006" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="171" birthdate="2008-01-01" gender="F" lastname="Liebhold" firstname="Lotta" license="0">
              <RESULTS>
                <RESULT resultid="698" eventid="1" swimtime="00:00:57.91" lane="1" heatid="1009" />
                <RESULT resultid="743" eventid="7" swimtime="00:00:24.18" lane="6" heatid="7002" />
                <RESULT resultid="721" eventid="11" swimtime="00:02:08.97" lane="4" heatid="11008">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:02.66" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="720" eventid="15" swimtime="00:20:21.78" lane="3" heatid="15001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:12.46" />
                    <SPLIT distance="200" swimtime="00:02:34.07" />
                    <SPLIT distance="300" swimtime="00:03:56.40" />
                    <SPLIT distance="400" swimtime="00:05:18.87" />
                    <SPLIT distance="500" swimtime="00:06:39.67" />
                    <SPLIT distance="600" swimtime="00:08:01.58" />
                    <SPLIT distance="700" swimtime="00:09:24.23" />
                    <SPLIT distance="800" swimtime="00:10:47.20" />
                    <SPLIT distance="900" swimtime="00:12:13.20" />
                    <SPLIT distance="1000" swimtime="00:13:40.24" />
                    <SPLIT distance="1100" swimtime="00:15:03.99" />
                    <SPLIT distance="1200" swimtime="00:16:29.37" />
                    <SPLIT distance="1300" swimtime="00:17:53.80" />
                    <SPLIT distance="1400" swimtime="00:19:14.28" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="749" eventid="16" swimtime="00:00:25.40" lane="1" heatid="16009" />
                <RESULT resultid="767" eventid="20" swimtime="00:09:54.00" lane="6" heatid="20002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:06.71" />
                    <SPLIT distance="200" swimtime="00:02:23.00" />
                    <SPLIT distance="300" swimtime="00:03:41.26" />
                    <SPLIT distance="400" swimtime="00:04:59.77" />
                    <SPLIT distance="500" swimtime="00:06:16.72" />
                    <SPLIT distance="600" swimtime="00:07:34.10" />
                    <SPLIT distance="700" swimtime="00:08:46.59" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="712" eventid="21" swimtime="00:01:00.11" lane="6" heatid="21003" />
                <RESULT resultid="731" eventid="25" swimtime="00:04:38.12" lane="8" heatid="25006">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:05.45" />
                    <SPLIT distance="200" swimtime="00:02:18.03" />
                    <SPLIT distance="300" swimtime="00:03:30.89" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="172" birthdate="2006-01-01" gender="F" lastname="Hollatz" firstname="Ronja" license="0">
              <RESULTS>
                <RESULT resultid="699" eventid="1" swimtime="00:00:57.83" lane="4" heatid="1008" />
                <RESULT resultid="742" eventid="7" swimtime="00:00:23.37" lane="3" heatid="7002" />
                <RESULT resultid="750" eventid="16" swimtime="00:00:25.55" lane="3" heatid="16008" />
                <RESULT resultid="711" eventid="21" swimtime="00:00:57.34" lane="8" heatid="21004" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="173" birthdate="2009-01-01" gender="F" lastname="Weber" firstname="Augusta Swantje" license="0">
              <RESULTS>
                <RESULT resultid="700" eventid="1" status="DNS" swimtime="00:00:00.00" lane="2" heatid="1007" />
                <RESULT resultid="722" eventid="11" status="DNS" swimtime="00:00:00.00" lane="6" heatid="11007" />
                <RESULT resultid="751" eventid="16" status="DNS" swimtime="00:00:00.00" lane="5" heatid="16006" />
                <RESULT resultid="713" eventid="21" status="DNS" swimtime="00:00:00.00" lane="8" heatid="21003" />
                <RESULT resultid="732" eventid="25" status="DNS" swimtime="00:00:00.00" lane="1" heatid="25005" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="174" birthdate="2010-01-01" gender="F" lastname="Rückert" firstname="Alma" license="0">
              <RESULTS>
                <RESULT resultid="701" eventid="1" swimtime="00:01:03.01" lane="6" heatid="1006" />
                <RESULT resultid="762" eventid="9" swimtime="00:00:28.54" lane="3" heatid="9002" />
                <RESULT resultid="723" eventid="11" swimtime="00:02:23.23" lane="1" heatid="11006">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:08.96" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="752" eventid="16" swimtime="00:00:27.95" lane="1" heatid="16006" />
                <RESULT resultid="714" eventid="21" swimtime="00:01:07.02" lane="5" heatid="21002" />
                <RESULT resultid="733" eventid="25" swimtime="00:05:10.33" lane="7" heatid="25004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:11.21" />
                    <SPLIT distance="200" swimtime="00:02:34.77" />
                    <SPLIT distance="300" swimtime="00:03:58.92" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="175" birthdate="2012-01-01" gender="F" lastname="Uhlig" firstname="Maike" license="0">
              <RESULTS>
                <RESULT resultid="702" eventid="1" swimtime="00:01:08.91" lane="2" heatid="1004" />
                <RESULT resultid="724" eventid="11" swimtime="00:02:38.63" lane="3" heatid="11004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:15.82" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="754" eventid="16" swimtime="00:00:30.71" lane="5" heatid="16003" />
                <RESULT resultid="735" eventid="25" swimtime="00:05:37.76" lane="6" heatid="25002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:17.78" />
                    <SPLIT distance="200" swimtime="00:02:46.23" />
                    <SPLIT distance="300" swimtime="00:04:15.08" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="176" birthdate="2010-01-01" gender="F" lastname="Hoffmann" firstname="Lydia" license="0">
              <RESULTS>
                <RESULT resultid="703" eventid="1" swimtime="00:01:08.33" lane="7" heatid="1004" />
                <RESULT resultid="763" eventid="9" swimtime="00:00:30.86" lane="4" heatid="9001" />
                <RESULT resultid="725" eventid="11" swimtime="00:02:37.73" lane="1" heatid="11004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:13.88" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="753" eventid="16" swimtime="00:00:29.90" lane="1" heatid="16004" />
                <RESULT resultid="765" eventid="20" swimtime="00:11:17.97" lane="4" heatid="20001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:13.13" />
                    <SPLIT distance="200" swimtime="00:02:41.73" />
                    <SPLIT distance="300" swimtime="00:04:11.79" />
                    <SPLIT distance="400" swimtime="00:05:41.04" />
                    <SPLIT distance="500" swimtime="00:07:07.04" />
                    <SPLIT distance="600" swimtime="00:08:35.29" />
                    <SPLIT distance="700" swimtime="00:10:02.02" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="715" eventid="21" swimtime="00:01:15.71" lane="7" heatid="21002" />
                <RESULT resultid="734" eventid="25" swimtime="00:05:40.74" lane="6" heatid="25003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:15.42" />
                    <SPLIT distance="200" swimtime="00:02:47.84" />
                    <SPLIT distance="300" swimtime="00:04:17.28" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="177" birthdate="2011-01-01" gender="F" lastname="Wirsching" firstname="Ellen" license="0">
              <RESULTS>
                <RESULT resultid="704" eventid="1" swimtime="00:01:16.78" lane="6" heatid="1003" />
                <RESULT resultid="726" eventid="11" swimtime="00:02:51.20" lane="4" heatid="11002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:22.10" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="755" eventid="16" swimtime="00:00:33.18" lane="6" heatid="16003" />
                <RESULT resultid="736" eventid="25" swimtime="00:05:58.84" lane="2" heatid="25002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:22.91" />
                    <SPLIT distance="200" swimtime="00:02:58.05" />
                    <SPLIT distance="300" swimtime="00:04:31.33" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="178" birthdate="2014-01-01" gender="F" lastname="Uhlig" firstname="Anna" license="0">
              <RESULTS>
                <RESULT resultid="705" eventid="1" swimtime="00:01:34.53" lane="7" heatid="1002" />
                <RESULT resultid="756" eventid="16" swimtime="00:00:42.50" lane="3" heatid="16001" />
                <RESULT resultid="746" eventid="23" swimtime="00:00:44.17" lane="4" heatid="23002" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="179" birthdate="2001-01-01" gender="M" lastname="Pohl" firstname="Enrico" license="0">
              <RESULTS>
                <RESULT resultid="706" eventid="2" swimtime="00:00:37.71" lane="3" heatid="2008" />
                <RESULT resultid="744" eventid="8" swimtime="00:00:15.62" lane="3" heatid="8004" />
                <RESULT resultid="727" eventid="12" swimtime="00:01:35.68" lane="1" heatid="12007">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:43.88" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="757" eventid="17" swimtime="00:00:17.33" lane="5" heatid="17008" />
                <RESULT resultid="716" eventid="22" swimtime="00:00:38.82" lane="3" heatid="22004" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="180" birthdate="2007-01-01" gender="M" lastname="Stuwe" firstname="Paul" license="0">
              <RESULTS>
                <RESULT resultid="707" eventid="2" swimtime="00:00:51.38" lane="3" heatid="2005" />
                <RESULT resultid="740" eventid="6" status="DSQ" swimtime="00:00:00.00" lane="8" heatid="6002" comment="Gesicht aus dem Wasser (Aufgegeben) nach 230 m">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:57.76" />
                    <SPLIT distance="200" swimtime="00:02:01.70" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="745" eventid="8" swimtime="00:00:20.35" lane="7" heatid="8002" />
                <RESULT resultid="719" eventid="15" swimtime="00:18:15.56" lane="7" heatid="15002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:04.89" />
                    <SPLIT distance="200" swimtime="00:02:17.69" />
                    <SPLIT distance="300" swimtime="00:03:30.52" />
                    <SPLIT distance="400" swimtime="00:04:43.76" />
                    <SPLIT distance="500" swimtime="00:05:56.87" />
                    <SPLIT distance="600" swimtime="00:07:10.64" />
                    <SPLIT distance="700" swimtime="00:08:25.03" />
                    <SPLIT distance="800" swimtime="00:09:37.85" />
                    <SPLIT distance="900" swimtime="00:10:52.23" />
                    <SPLIT distance="1000" swimtime="00:12:06.90" />
                    <SPLIT distance="1100" swimtime="00:13:22.30" />
                    <SPLIT distance="1200" swimtime="00:14:36.82" />
                    <SPLIT distance="1300" swimtime="00:15:52.16" />
                    <SPLIT distance="1400" swimtime="00:17:04.26" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="758" eventid="17" swimtime="00:00:22.87" lane="7" heatid="17006" />
                <RESULT resultid="766" eventid="20" swimtime="00:08:50.03" lane="5" heatid="20003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:59.82" />
                    <SPLIT distance="200" swimtime="00:02:05.21" />
                    <SPLIT distance="300" swimtime="00:03:11.25" />
                    <SPLIT distance="400" swimtime="00:04:18.36" />
                    <SPLIT distance="500" swimtime="00:05:26.56" />
                    <SPLIT distance="600" swimtime="00:06:36.20" />
                    <SPLIT distance="700" swimtime="00:07:44.21" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="717" eventid="22" swimtime="00:00:48.39" lane="7" heatid="22003" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="181" birthdate="2011-01-01" gender="M" lastname="Knöfel" firstname="Florian" license="0">
              <RESULTS>
                <RESULT resultid="708" eventid="2" swimtime="00:01:15.13" lane="6" heatid="2003" />
                <RESULT resultid="764" eventid="10" swimtime="00:00:33.74" lane="5" heatid="10001" />
                <RESULT resultid="729" eventid="12" swimtime="00:02:49.90" lane="1" heatid="12003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:24.23" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="759" eventid="17" swimtime="00:00:31.73" lane="5" heatid="17003" />
                <RESULT resultid="718" eventid="22" swimtime="00:01:18.68" lane="7" heatid="22001" />
                <RESULT resultid="738" eventid="26" swimtime="00:06:05.12" lane="7" heatid="26002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:30.42" />
                    <SPLIT distance="200" swimtime="00:03:04.70" />
                    <SPLIT distance="300" swimtime="00:04:37.64" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="182" birthdate="2011-01-01" gender="M" lastname="Bartels" firstname="Constantin" license="0">
              <RESULTS>
                <RESULT resultid="709" eventid="2" swimtime="00:01:28.39" lane="3" heatid="2002" />
                <RESULT resultid="730" eventid="12" swimtime="00:03:15.35" lane="4" heatid="12002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:31.99" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="760" eventid="17" swimtime="00:00:41.36" lane="3" heatid="17002" />
                <RESULT resultid="739" eventid="26" swimtime="00:06:48.72" lane="1" heatid="26002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:35.85" />
                    <SPLIT distance="200" swimtime="00:03:21.50" />
                    <SPLIT distance="300" swimtime="00:05:07.16" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="183" birthdate="2016-01-01" gender="M" lastname="Stuwe" firstname="Piet" license="0">
              <RESULTS>
                <RESULT resultid="761" eventid="17" swimtime="00:00:47.49" lane="5" heatid="17001" />
                <RESULT resultid="747" eventid="24" status="DSQ" swimtime="00:00:52.36" lane="1" heatid="24001" comment="falscher Schwimmstil (Beinwechselschlag) bei 15m" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="233" birthdate="1998-01-01" gender="M" lastname="Rose" firstname="Jonas" license="0">
              <RESULTS>
                <RESULT resultid="978" eventid="6" status="DNS" swimtime="00:00:00.00" lane="7" heatid="6002" />
                <RESULT resultid="979" eventid="15" status="DNS" swimtime="00:00:00.00" lane="4" heatid="15002" />
                <RESULT resultid="980" eventid="20" status="DNS" swimtime="00:00:00.00" lane="4" heatid="20003" />
                <RESULT resultid="981" eventid="22" status="DNS" swimtime="00:00:00.00" lane="7" heatid="22004" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY number="1" gender="X" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="969" eventid="13" swimtime="00:01:25.74" lane="3" heatid="13003">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="179" number="1" />
                    <RELAYPOSITION athleteid="170" number="2" />
                    <RELAYPOSITION athleteid="180" number="3" />
                    <RELAYPOSITION athleteid="171" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="2" gender="X" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="970" eventid="13" swimtime="00:02:12.60" lane="7" heatid="13002">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="174" number="1" />
                    <RELAYPOSITION athleteid="181" number="2" />
                    <RELAYPOSITION athleteid="176" number="3" />
                    <RELAYPOSITION athleteid="182" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
      </CLUBS>
    </MEET>
  </MEETS>
</LENEX>
