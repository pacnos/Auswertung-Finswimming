<?xml version="1.0" encoding="UTF-8"?>
<LENEX version="3.0">
  <CONSTRUCTOR name="EasyWk" version="5.24 BETA" registration="">
    <CONTACT name="Bjoern Stickan" internet="http://www.easywk.de" email="info@easywk.de" />
  </CONSTRUCTOR>
  <MEETS>
    <MEET city="Dresden" course="LCM" name="Sparkassen Landesjugendspiele 2023 Zeig Dein Sporttalent!" nation="GER" organizer="Sächsischer Schwimm-Verband e.V. / Dresdner Delphine e.V." hostclub="Landessportbund Sachsen e.V." deadline="2023-06-23" timing="AUTOMATIC">
      <CONTACT city="Leipzig" email="landesjugendspiele2023@egd-tb.info" fax="+49-341-4426911" internet="https://dsvdaten.dsv.de/File.aspx?F=WKInfo&amp;File=1792023.pdf" name="Brandenburg, Thilo" phone="+49-178-8150839" street="Zum Leutzscher Holz 26" zip="04178" />
      <AGEDATE type="YEAR" value="2023-01-01" />
      <SESSIONS>
        <SESSION number="1" date="2023-07-01" daytime="10:00" officialmeeting="09:30" warmupfrom="09:00">
          <EVENTS>
            <EVENT eventid="1" number="1" gender="F" round="TIM">
              <SWIMSTYLE stroke="MEDLEY" relaycount="1" distance="200" />
              <HEATS>
                <HEAT heatid="1001" number="1" />
                <HEAT heatid="1002" number="2" />
                <HEAT heatid="1003" number="3" />
                <HEAT heatid="1004" number="4" />
                <HEAT heatid="1005" number="5" />
                <HEAT heatid="1006" number="6" />
                <HEAT heatid="1007" number="7" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="10" agemin="10" name="Jahrgang 2013">
                  <RANKINGS>
                    <RANKING place="1" resultid="7" />
                    <RANKING place="4" resultid="846" />
                    <RANKING place="5" resultid="5188" />
                    <RANKING place="2" resultid="5438" />
                    <RANKING place="3" resultid="5572" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2" agemax="11" agemin="11" name="Jahrgang 2012">
                  <RANKINGS>
                    <RANKING place="5" resultid="14" />
                    <RANKING place="6" resultid="2127" />
                    <RANKING place="3" resultid="4736" />
                    <RANKING place="7" resultid="5228" />
                    <RANKING place="2" resultid="5339" />
                    <RANKING place="9" resultid="5668" />
                    <RANKING place="4" resultid="5709" />
                    <RANKING place="8" resultid="6033" />
                    <RANKING place="1" resultid="6062" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="13" agemin="12" name="Jahrgang 2010/2011">
                  <RANKINGS>
                    <RANKING place="7" resultid="145" />
                    <RANKING place="6" resultid="153" />
                    <RANKING place="4" resultid="978" />
                    <RANKING place="11" resultid="1948" />
                    <RANKING place="16" resultid="2064" />
                    <RANKING place="2" resultid="2143" />
                    <RANKING place="17" resultid="4028" />
                    <RANKING place="9" resultid="4059" />
                    <RANKING place="18" resultid="4544" />
                    <RANKING place="13" resultid="4926" />
                    <RANKING place="5" resultid="5236" />
                    <RANKING place="14" resultid="5326" />
                    <RANKING place="19" resultid="5365" />
                    <RANKING place="8" resultid="5400" />
                    <RANKING place="3" resultid="5435" />
                    <RANKING place="15" resultid="5460" />
                    <RANKING place="12" resultid="5556" />
                    <RANKING place="21" resultid="5604" />
                    <RANKING place="20" resultid="5704" />
                    <RANKING place="10" resultid="5798" />
                    <RANKING place="1" resultid="6135" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6" agemax="15" agemin="14" name="Jahrgang 2008/2009">
                  <RANKINGS>
                    <RANKING place="11" resultid="3724" />
                    <RANKING place="1" resultid="4577" />
                    <RANKING place="4" resultid="4992" />
                    <RANKING place="2" resultid="5351" />
                    <RANKING place="5" resultid="5496" />
                    <RANKING place="7" resultid="5608" />
                    <RANKING place="10" resultid="5663" />
                    <RANKING place="8" resultid="5872" />
                    <RANKING place="6" resultid="5961" />
                    <RANKING place="9" resultid="6138" />
                    <RANKING place="3" resultid="6273" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8" agemax="17" agemin="16" name="Jahrgang 2006/2007">
                  <RANKINGS>
                    <RANKING place="4" resultid="1912" />
                    <RANKING place="3" resultid="4647" />
                    <RANKING place="1" resultid="4671" />
                    <RANKING place="2" resultid="6349" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="2" number="2" gender="M" round="TIM">
              <SWIMSTYLE stroke="MEDLEY" relaycount="1" distance="200" />
              <HEATS>
                <HEAT heatid="2001" number="1" />
                <HEAT heatid="2002" number="2" />
                <HEAT heatid="2003" number="3" />
                <HEAT heatid="2004" number="4" />
                <HEAT heatid="2005" number="5" />
                <HEAT heatid="2006" number="6" />
                <HEAT heatid="2007" number="7" />
                <HEAT heatid="2008" number="8" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="10" agemin="10" name="Jahrgang 2013">
                  <RANKINGS>
                    <RANKING place="1" resultid="831" />
                    <RANKING place="10" resultid="4173" />
                    <RANKING place="7" resultid="4774" />
                    <RANKING place="5" resultid="5258" />
                    <RANKING place="9" resultid="5335" />
                    <RANKING place="8" resultid="5536" />
                    <RANKING place="2" resultid="5623" />
                    <RANKING place="4" resultid="5885" />
                    <RANKING place="3" resultid="5949" />
                    <RANKING place="6" resultid="6258" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2" agemax="11" agemin="11" name="Jahrgang 2012">
                  <RANKINGS>
                    <RANKING place="1" resultid="121" />
                    <RANKING place="2" resultid="185" />
                    <RANKING place="5" resultid="824" />
                    <RANKING place="11" resultid="995" />
                    <RANKING place="4" resultid="2109" />
                    <RANKING place="12" resultid="4063" />
                    <RANKING place="3" resultid="4722" />
                    <RANKING place="7" resultid="5515" />
                    <RANKING place="13" resultid="5564" />
                    <RANKING place="8" resultid="5684" />
                    <RANKING place="6" resultid="5814" />
                    <RANKING place="10" resultid="5937" />
                    <RANKING place="9" resultid="6291" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="13" agemin="12" name="Jahrgang 2010/2011">
                  <RANKINGS>
                    <RANKING place="7" resultid="113" />
                    <RANKING place="6" resultid="137" />
                    <RANKING place="4" resultid="796" />
                    <RANKING place="3" resultid="875" />
                    <RANKING place="19" resultid="1934" />
                    <RANKING place="17" resultid="2025" />
                    <RANKING place="11" resultid="4020" />
                    <RANKING place="13" resultid="4075" />
                    <RANKING place="12" resultid="4589" />
                    <RANKING place="15" resultid="5270" />
                    <RANKING place="20" resultid="5282" />
                    <RANKING place="9" resultid="5423" />
                    <RANKING place="16" resultid="5658" />
                    <RANKING place="5" resultid="5697" />
                    <RANKING place="18" resultid="5738" />
                    <RANKING place="8" resultid="5745" />
                    <RANKING place="14" resultid="5879" />
                    <RANKING place="21" resultid="5894" />
                    <RANKING place="1" resultid="5923" />
                    <RANKING place="2" resultid="6220" />
                    <RANKING place="10" resultid="6326" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6" agemax="15" agemin="14" name="Jahrgang 2008/2009">
                  <RANKINGS>
                    <RANKING place="3" resultid="3716" />
                    <RANKING place="4" resultid="3836" />
                    <RANKING place="2" resultid="5384" />
                    <RANKING place="1" resultid="5900" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8" agemax="17" agemin="16" name="Jahrgang 2006/2007">
                  <RANKINGS>
                    <RANKING place="4" resultid="3488" />
                    <RANKING place="5" resultid="4573" />
                    <RANKING place="1" resultid="4706" />
                    <RANKING place="3" resultid="5131" />
                    <RANKING place="2" resultid="5313" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="39" number="101" gender="F" round="TIM">
              <SWIMSTYLE stroke="SURFACE" name="200 Flossenschwimmen Frauen" relaycount="1" distance="200" />
              <HEATS>
                <HEAT heatid="39001" number="1" />
                <HEAT heatid="39002" number="2" />
                <HEAT heatid="39003" number="3" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="9" agemin="8" name="Jahrgang 2014/2015">
                  <RANKINGS>
                    <RANKING place="2" resultid="33" />
                    <RANKING place="1" resultid="41" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2" agemax="11" agemin="10" name="Jahrgang 2012/2013">
                  <RANKINGS>
                    <RANKING place="4" resultid="579" />
                    <RANKING place="2" resultid="1532" />
                    <RANKING place="1" resultid="1564" />
                    <RANKING place="3" resultid="1568" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3" agemax="14" agemin="12" name="Jahrgang 2009 bis 2011">
                  <RANKINGS>
                    <RANKING place="6" resultid="25" />
                    <RANKING place="2" resultid="29" />
                    <RANKING place="9" resultid="573" />
                    <RANKING place="7" resultid="599" />
                    <RANKING place="8" resultid="1546" />
                    <RANKING place="3" resultid="1582" />
                    <RANKING place="5" resultid="2153" />
                    <RANKING place="4" resultid="2182" />
                    <RANKING place="1" resultid="4180" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="17" agemin="15" name="Jahrgang 2006 bis 2008">
                  <RANKINGS>
                    <RANKING place="4" resultid="583" />
                    <RANKING place="6" resultid="595" />
                    <RANKING place="2" resultid="1535" />
                    <RANKING place="1" resultid="2176" />
                    <RANKING place="3" resultid="3997" />
                    <RANKING place="5" resultid="4001" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="40" number="102" gender="M" round="TIM">
              <SWIMSTYLE stroke="SURFACE" name="200 Flossenschwimmen Männer" relaycount="1" distance="200" />
              <HEATS>
                <HEAT heatid="40001" number="1" />
                <HEAT heatid="40002" number="2" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="9" agemin="8" name="Jahrgang 2014/2015">
                  <RANKINGS>
                    <RANKING place="3" resultid="37" />
                    <RANKING place="2" resultid="45" />
                    <RANKING place="1" resultid="587" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2" agemax="11" agemin="10" name="Jahrgang 2012/2013">
                  <RANKINGS>
                    <RANKING place="6" resultid="565" />
                    <RANKING place="3" resultid="569" />
                    <RANKING place="2" resultid="591" />
                    <RANKING place="5" resultid="606" />
                    <RANKING place="1" resultid="1542" />
                    <RANKING place="4" resultid="2156" />
                    <RANKING place="7" resultid="2189" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3" agemax="14" agemin="12" name="Jahrgang 2009 bis 2011">
                  <RANKINGS>
                    <RANKING place="1" resultid="2148" />
                    <RANKING place="3" resultid="2159" />
                    <RANKING place="2" resultid="2193" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="17" agemin="15" name="Jahrgang 2006 bis 2008">
                  <RANKINGS>
                    <RANKING place="1" resultid="603" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="3" number="3" gender="F" round="TIM">
              <SWIMSTYLE stroke="BREAST" relaycount="1" distance="100" />
              <HEATS>
                <HEAT heatid="3001" number="1" />
                <HEAT heatid="3002" number="2" />
                <HEAT heatid="3003" number="3" />
                <HEAT heatid="3004" number="4" />
                <HEAT heatid="3005" number="5" />
                <HEAT heatid="3006" number="6" />
                <HEAT heatid="3007" number="7" />
                <HEAT heatid="3008" number="8" />
                <HEAT heatid="3009" number="9" />
                <HEAT heatid="3010" number="10" />
                <HEAT heatid="3011" number="11" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="10" agemin="10" name="Jahrgang 2013">
                  <RANKINGS>
                    <RANKING place="5" resultid="470" />
                    <RANKING place="2" resultid="898" />
                    <RANKING place="8" resultid="3828" />
                    <RANKING place="17" resultid="4125" />
                    <RANKING place="16" resultid="4157" />
                    <RANKING place="14" resultid="4256" />
                    <RANKING place="12" resultid="4259" />
                    <RANKING place="10" resultid="4613" />
                    <RANKING place="13" resultid="4632" />
                    <RANKING place="3" resultid="4746" />
                    <RANKING place="18" resultid="4956" />
                    <RANKING place="7" resultid="5094" />
                    <RANKING place="11" resultid="5161" />
                    <RANKING place="1" resultid="5217" />
                    <RANKING place="6" resultid="5475" />
                    <RANKING place="15" resultid="5778" />
                    <RANKING place="4" resultid="5827" />
                    <RANKING place="9" resultid="6047" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2" agemax="11" agemin="11" name="Jahrgang 2012">
                  <RANKINGS>
                    <RANKING place="6" resultid="177" />
                    <RANKING place="5" resultid="961" />
                    <RANKING place="9" resultid="1600" />
                    <RANKING place="19" resultid="1648" />
                    <RANKING place="12" resultid="2116" />
                    <RANKING place="8" resultid="2126" />
                    <RANKING place="10" resultid="4810" />
                    <RANKING place="18" resultid="4870" />
                    <RANKING place="15" resultid="5033" />
                    <RANKING place="1" resultid="5340" />
                    <RANKING place="17" resultid="5490" />
                    <RANKING place="21" resultid="5615" />
                    <RANKING place="2" resultid="5635" />
                    <RANKING place="7" resultid="5642" />
                    <RANKING place="20" resultid="5669" />
                    <RANKING place="14" resultid="5717" />
                    <RANKING place="13" resultid="5929" />
                    <RANKING place="16" resultid="6021" />
                    <RANKING place="11" resultid="6175" />
                    <RANKING place="4" resultid="6232" />
                    <RANKING place="3" resultid="6315" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="13" agemin="12" name="Jahrgang 2010/2011">
                  <RANKINGS>
                    <RANKING place="4" resultid="129" />
                    <RANKING place="9" resultid="146" />
                    <RANKING place="6" resultid="169" />
                    <RANKING place="1" resultid="234" />
                    <RANKING place="3" resultid="611" />
                    <RANKING place="2" resultid="3454" />
                    <RANKING place="12" resultid="4029" />
                    <RANKING place="19" resultid="4107" />
                    <RANKING place="29" resultid="4131" />
                    <RANKING place="17" resultid="4545" />
                    <RANKING place="22" resultid="4694" />
                    <RANKING place="21" resultid="4863" />
                    <RANKING place="7" resultid="4877" />
                    <RANKING place="23" resultid="4999" />
                    <RANKING place="25" resultid="5082" />
                    <RANKING place="14" resultid="5145" />
                    <RANKING place="11" resultid="5205" />
                    <RANKING place="8" resultid="5255" />
                    <RANKING place="18" resultid="5278" />
                    <RANKING place="27" resultid="5366" />
                    <RANKING place="5" resultid="5389" />
                    <RANKING place="10" resultid="5401" />
                    <RANKING place="24" resultid="5758" />
                    <RANKING place="15" resultid="5773" />
                    <RANKING place="28" resultid="5784" />
                    <RANKING place="20" resultid="5787" />
                    <RANKING place="26" resultid="6002" />
                    <RANKING place="30" resultid="6077" />
                    <RANKING place="16" resultid="6281" />
                    <RANKING place="13" resultid="6359" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6" agemax="15" agemin="14" name="Jahrgang 2008/2009">
                  <RANKINGS>
                    <RANKING place="1" resultid="3823" />
                    <RANKING place="2" resultid="4884" />
                    <RANKING place="6" resultid="5319" />
                    <RANKING place="3" resultid="5649" />
                    <RANKING place="4" resultid="5917" />
                    <RANKING place="5" resultid="6187" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8" agemax="17" agemin="16" name="Jahrgang 2006/2007">
                  <RANKINGS>
                    <RANKING place="2" resultid="4621" />
                    <RANKING place="1" resultid="4700" />
                    <RANKING place="3" resultid="4837" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="4" number="4" gender="M" round="TIM">
              <SWIMSTYLE stroke="BREAST" relaycount="1" distance="100" />
              <HEATS>
                <HEAT heatid="4001" number="1" />
                <HEAT heatid="4002" number="2" />
                <HEAT heatid="4003" number="3" />
                <HEAT heatid="4004" number="4" />
                <HEAT heatid="4005" number="5" />
                <HEAT heatid="4006" number="6" />
                <HEAT heatid="4007" number="7" />
                <HEAT heatid="4008" number="8" />
                <HEAT heatid="4009" number="9" />
                <HEAT heatid="4010" number="10" />
                <HEAT heatid="4011" number="11" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="10" agemin="10" name="Jahrgang 2013">
                  <RANKINGS>
                    <RANKING place="4" resultid="853" />
                    <RANKING place="9" resultid="1627" />
                    <RANKING place="2" resultid="1633" />
                    <RANKING place="3" resultid="4038" />
                    <RANKING place="8" resultid="4097" />
                    <RANKING place="7" resultid="4757" />
                    <RANKING place="11" resultid="4775" />
                    <RANKING place="12" resultid="4981" />
                    <RANKING place="10" resultid="5061" />
                    <RANKING place="1" resultid="5584" />
                    <RANKING place="5" resultid="5950" />
                    <RANKING place="13" resultid="6124" />
                    <RANKING place="6" resultid="6196" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2" agemax="11" agemin="11" name="Jahrgang 2012">
                  <RANKINGS>
                    <RANKING place="13" resultid="161" />
                    <RANKING place="3" resultid="823" />
                    <RANKING place="17" resultid="860" />
                    <RANKING place="10" resultid="2120" />
                    <RANKING place="1" resultid="3459" />
                    <RANKING place="16" resultid="3751" />
                    <RANKING place="11" resultid="4064" />
                    <RANKING place="20" resultid="4167" />
                    <RANKING place="12" resultid="4240" />
                    <RANKING place="14" resultid="4716" />
                    <RANKING place="6" resultid="4795" />
                    <RANKING place="9" resultid="4824" />
                    <RANKING place="4" resultid="5167" />
                    <RANKING place="5" resultid="5305" />
                    <RANKING place="8" resultid="5523" />
                    <RANKING place="18" resultid="5546" />
                    <RANKING place="19" resultid="5807" />
                    <RANKING place="2" resultid="5815" />
                    <RANKING place="15" resultid="5848" />
                    <RANKING place="7" resultid="6099" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="13" agemin="12" name="Jahrgang 2010/2011">
                  <RANKINGS>
                    <RANKING place="6" resultid="138" />
                    <RANKING place="1" resultid="240" />
                    <RANKING place="3" resultid="773" />
                    <RANKING place="8" resultid="1962" />
                    <RANKING place="4" resultid="3445" />
                    <RANKING place="19" resultid="3815" />
                    <RANKING place="24" resultid="3850" />
                    <RANKING place="9" resultid="4283" />
                    <RANKING place="7" resultid="4464" />
                    <RANKING place="10" resultid="4551" />
                    <RANKING place="15" resultid="4567" />
                    <RANKING place="2" resultid="4625" />
                    <RANKING place="21" resultid="4638" />
                    <RANKING place="13" resultid="4890" />
                    <RANKING place="18" resultid="4897" />
                    <RANKING place="22" resultid="5262" />
                    <RANKING place="14" resultid="5271" />
                    <RANKING place="5" resultid="5451" />
                    <RANKING place="16" resultid="5739" />
                    <RANKING place="11" resultid="5742" />
                    <RANKING place="12" resultid="5880" />
                    <RANKING place="20" resultid="5895" />
                    <RANKING place="17" resultid="6029" />
                    <RANKING place="23" resultid="6209" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6" agemax="15" agemin="14" name="Jahrgang 2008/2009">
                  <RANKINGS>
                    <RANKING place="3" resultid="3778" />
                    <RANKING place="9" resultid="4103" />
                    <RANKING place="6" resultid="4314" />
                    <RANKING place="16" resultid="4536" />
                    <RANKING place="10" resultid="4596" />
                    <RANKING place="11" resultid="4659" />
                    <RANKING place="2" resultid="4781" />
                    <RANKING place="15" resultid="4804" />
                    <RANKING place="14" resultid="4817" />
                    <RANKING place="7" resultid="4849" />
                    <RANKING place="12" resultid="4903" />
                    <RANKING place="5" resultid="4949" />
                    <RANKING place="4" resultid="5359" />
                    <RANKING place="13" resultid="5681" />
                    <RANKING place="1" resultid="5835" />
                    <RANKING place="8" resultid="6080" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8" agemax="17" agemin="16" name="Jahrgang 2006/2007">
                  <RANKINGS>
                    <RANKING place="1" resultid="3469" />
                    <RANKING place="5" resultid="3799" />
                    <RANKING place="2" resultid="4293" />
                    <RANKING place="3" resultid="4831" />
                    <RANKING place="4" resultid="5580" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="5" number="5" gender="F" round="TIM">
              <SWIMSTYLE stroke="FLY" relaycount="1" distance="50" />
              <HEATS>
                <HEAT heatid="5001" number="1" />
                <HEAT heatid="5002" number="2" />
                <HEAT heatid="5003" number="3" />
                <HEAT heatid="5004" number="4" />
                <HEAT heatid="5005" number="5" />
                <HEAT heatid="5006" number="6" />
                <HEAT heatid="5007" number="7" />
                <HEAT heatid="5008" number="8" />
                <HEAT heatid="5009" number="9" />
                <HEAT heatid="5010" number="10" />
                <HEAT heatid="5011" number="11" />
                <HEAT heatid="5012" number="12" />
                <HEAT heatid="5013" number="13" />
                <HEAT heatid="5014" number="14" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="10" agemin="10" name="Jahrgang 2013">
                  <RANKINGS>
                    <RANKING place="1" resultid="8" />
                    <RANKING place="5" resultid="845" />
                    <RANKING place="3" resultid="891" />
                    <RANKING place="14" resultid="953" />
                    <RANKING place="7" resultid="2123" />
                    <RANKING place="13" resultid="4260" />
                    <RANKING place="9" resultid="4614" />
                    <RANKING place="11" resultid="4689" />
                    <RANKING place="15" resultid="4957" />
                    <RANKING place="10" resultid="5139" />
                    <RANKING place="12" resultid="5189" />
                    <RANKING place="6" resultid="5218" />
                    <RANKING place="4" resultid="5439" />
                    <RANKING place="8" resultid="5476" />
                    <RANKING place="2" resultid="5573" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2" agemax="11" agemin="11" name="Jahrgang 2012">
                  <RANKINGS>
                    <RANKING place="3" resultid="15" />
                    <RANKING place="15" resultid="178" />
                    <RANKING place="7" resultid="960" />
                    <RANKING place="13" resultid="1611" />
                    <RANKING place="10" resultid="1617" />
                    <RANKING place="21" resultid="1654" />
                    <RANKING place="6" resultid="1957" />
                    <RANKING place="8" resultid="4737" />
                    <RANKING place="28" resultid="4857" />
                    <RANKING place="26" resultid="4871" />
                    <RANKING place="20" resultid="4910" />
                    <RANKING place="17" resultid="4917" />
                    <RANKING place="25" resultid="5034" />
                    <RANKING place="24" resultid="5105" />
                    <RANKING place="11" resultid="5177" />
                    <RANKING place="9" resultid="5229" />
                    <RANKING place="2" resultid="5341" />
                    <RANKING place="5" resultid="5710" />
                    <RANKING place="23" resultid="5718" />
                    <RANKING place="27" resultid="5793" />
                    <RANKING place="4" resultid="5841" />
                    <RANKING place="18" resultid="5930" />
                    <RANKING place="22" resultid="5972" />
                    <RANKING place="29" resultid="6022" />
                    <RANKING place="12" resultid="6034" />
                    <RANKING place="1" resultid="6063" />
                    <RANKING place="19" resultid="6176" />
                    <RANKING place="14" resultid="6233" />
                    <RANKING place="16" resultid="6316" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="13" agemin="12" name="Jahrgang 2010/2011">
                  <RANKINGS>
                    <RANKING place="2" resultid="130" />
                    <RANKING place="9" resultid="154" />
                    <RANKING place="4" resultid="170" />
                    <RANKING place="16" resultid="977" />
                    <RANKING place="5" resultid="2142" />
                    <RANKING place="29" resultid="3743" />
                    <RANKING place="8" resultid="4060" />
                    <RANKING place="26" resultid="4556" />
                    <RANKING place="14" resultid="4864" />
                    <RANKING place="20" resultid="4927" />
                    <RANKING place="28" resultid="5000" />
                    <RANKING place="19" resultid="5083" />
                    <RANKING place="13" resultid="5206" />
                    <RANKING place="10" resultid="5237" />
                    <RANKING place="24" resultid="5279" />
                    <RANKING place="11" resultid="5327" />
                    <RANKING place="17" resultid="5367" />
                    <RANKING place="7" resultid="5390" />
                    <RANKING place="12" resultid="5402" />
                    <RANKING place="6" resultid="5436" />
                    <RANKING place="14" resultid="5461" />
                    <RANKING place="22" resultid="5605" />
                    <RANKING place="25" resultid="5705" />
                    <RANKING place="23" resultid="5774" />
                    <RANKING place="27" resultid="5785" />
                    <RANKING place="3" resultid="5799" />
                    <RANKING place="30" resultid="6003" />
                    <RANKING place="1" resultid="6136" />
                    <RANKING place="18" resultid="6282" />
                    <RANKING place="21" resultid="6362" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6" agemax="15" agemin="14" name="Jahrgang 2008/2009">
                  <RANKINGS>
                    <RANKING place="8" resultid="3474" />
                    <RANKING place="21" resultid="3723" />
                    <RANKING place="3" resultid="4578" />
                    <RANKING place="13" resultid="4742" />
                    <RANKING place="16" resultid="4885" />
                    <RANKING place="5" resultid="4940" />
                    <RANKING place="10" resultid="4993" />
                    <RANKING place="12" resultid="5058" />
                    <RANKING place="18" resultid="5320" />
                    <RANKING place="4" resultid="5352" />
                    <RANKING place="2" resultid="5431" />
                    <RANKING place="20" resultid="5454" />
                    <RANKING place="19" resultid="5664" />
                    <RANKING place="15" resultid="5873" />
                    <RANKING place="9" resultid="5913" />
                    <RANKING place="17" resultid="5918" />
                    <RANKING place="11" resultid="5962" />
                    <RANKING place="1" resultid="6041" />
                    <RANKING place="7" resultid="6139" />
                    <RANKING place="14" resultid="6156" />
                    <RANKING place="6" resultid="6274" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8" agemax="17" agemin="16" name="Jahrgang 2006/2007">
                  <RANKINGS>
                    <RANKING place="7" resultid="4648" />
                    <RANKING place="3" resultid="4672" />
                    <RANKING place="5" resultid="4701" />
                    <RANKING place="6" resultid="4729" />
                    <RANKING place="9" resultid="4838" />
                    <RANKING place="8" resultid="5010" />
                    <RANKING place="4" resultid="5486" />
                    <RANKING place="1" resultid="6160" />
                    <RANKING place="2" resultid="6350" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="6" number="6" gender="M" round="TIM">
              <SWIMSTYLE stroke="FLY" relaycount="1" distance="50" />
              <HEATS>
                <HEAT heatid="6001" number="1" />
                <HEAT heatid="6002" number="2" />
                <HEAT heatid="6003" number="3" />
                <HEAT heatid="6004" number="4" />
                <HEAT heatid="6005" number="5" />
                <HEAT heatid="6006" number="6" />
                <HEAT heatid="6007" number="7" />
                <HEAT heatid="6008" number="8" />
                <HEAT heatid="6009" number="9" />
                <HEAT heatid="6010" number="10" />
                <HEAT heatid="6011" number="11" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="10" agemin="10" name="Jahrgang 2013">
                  <RANKINGS>
                    <RANKING place="1" resultid="830" />
                    <RANKING place="3" resultid="946" />
                    <RANKING place="2" resultid="3439" />
                    <RANKING place="14" resultid="3804" />
                    <RANKING place="12" resultid="3807" />
                    <RANKING place="7" resultid="4050" />
                    <RANKING place="8" resultid="4174" />
                    <RANKING place="9" resultid="4246" />
                    <RANKING place="11" resultid="5336" />
                    <RANKING place="10" resultid="5537" />
                    <RANKING place="4" resultid="5624" />
                    <RANKING place="5" resultid="5886" />
                    <RANKING place="13" resultid="6125" />
                    <RANKING place="6" resultid="6259" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2" agemax="11" agemin="11" name="Jahrgang 2012">
                  <RANKINGS>
                    <RANKING place="3" resultid="122" />
                    <RANKING place="2" resultid="186" />
                    <RANKING place="20" resultid="816" />
                    <RANKING place="9" resultid="918" />
                    <RANKING place="13" resultid="994" />
                    <RANKING place="18" resultid="1002" />
                    <RANKING place="5" resultid="2108" />
                    <RANKING place="21" resultid="2112" />
                    <RANKING place="14" resultid="2119" />
                    <RANKING place="12" resultid="4241" />
                    <RANKING place="17" resultid="4266" />
                    <RANKING place="4" resultid="4723" />
                    <RANKING place="19" resultid="4825" />
                    <RANKING place="6" resultid="5168" />
                    <RANKING place="11" resultid="5412" />
                    <RANKING place="8" resultid="5516" />
                    <RANKING place="16" resultid="5565" />
                    <RANKING place="7" resultid="5685" />
                    <RANKING place="10" resultid="5938" />
                    <RANKING place="1" resultid="6183" />
                    <RANKING place="15" resultid="6292" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="13" agemin="12" name="Jahrgang 2010/2011">
                  <RANKINGS>
                    <RANKING place="3" resultid="114" />
                    <RANKING place="6" resultid="795" />
                    <RANKING place="1" resultid="874" />
                    <RANKING place="12" resultid="3477" />
                    <RANKING place="7" resultid="4021" />
                    <RANKING place="11" resultid="4284" />
                    <RANKING place="5" resultid="4465" />
                    <RANKING place="22" resultid="4539" />
                    <RANKING place="8" resultid="4590" />
                    <RANKING place="15" resultid="4603" />
                    <RANKING place="18" resultid="4608" />
                    <RANKING place="2" resultid="4626" />
                    <RANKING place="20" resultid="4891" />
                    <RANKING place="21" resultid="5263" />
                    <RANKING place="13" resultid="5272" />
                    <RANKING place="17" resultid="5283" />
                    <RANKING place="9" resultid="5452" />
                    <RANKING place="14" resultid="5659" />
                    <RANKING place="10" resultid="5746" />
                    <RANKING place="19" resultid="5896" />
                    <RANKING place="4" resultid="5924" />
                    <RANKING place="16" resultid="6327" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6" agemax="15" agemin="14" name="Jahrgang 2008/2009">
                  <RANKINGS>
                    <RANKING place="16" resultid="3771" />
                    <RANKING place="11" resultid="3777" />
                    <RANKING place="2" resultid="4104" />
                    <RANKING place="8" resultid="4315" />
                    <RANKING place="7" resultid="4660" />
                    <RANKING place="6" resultid="4782" />
                    <RANKING place="14" resultid="4818" />
                    <RANKING place="3" resultid="4850" />
                    <RANKING place="13" resultid="4904" />
                    <RANKING place="5" resultid="4950" />
                    <RANKING place="4" resultid="5360" />
                    <RANKING place="10" resultid="5385" />
                    <RANKING place="15" resultid="5428" />
                    <RANKING place="9" resultid="5998" />
                    <RANKING place="1" resultid="6017" />
                    <RANKING place="12" resultid="6095" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8" agemax="17" agemin="16" name="Jahrgang 2006/2007">
                  <RANKINGS>
                    <RANKING place="3" resultid="3468" />
                    <RANKING place="5" resultid="3487" />
                    <RANKING place="7" resultid="4294" />
                    <RANKING place="4" resultid="4574" />
                    <RANKING place="1" resultid="4707" />
                    <RANKING place="6" resultid="4832" />
                    <RANKING place="2" resultid="5132" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="41" number="103" gender="F" round="TIM">
              <SWIMSTYLE stroke="APNEA" name="25 Apnoe Frauen" relaycount="1" distance="25" />
              <HEATS>
                <HEAT heatid="41001" number="1" />
                <HEAT heatid="41002" number="2" />
                <HEAT heatid="41003" number="3" />
                <HEAT heatid="41004" number="4" />
                <HEAT heatid="41005" number="5" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="2" agemax="11" agemin="10" name="Jahrgang 2012/2013">
                  <RANKINGS>
                    <RANKING place="2" resultid="580" />
                    <RANKING place="5" resultid="1531" />
                    <RANKING place="1" resultid="1563" />
                    <RANKING place="6" resultid="1567" />
                    <RANKING place="3" resultid="1576" />
                    <RANKING place="4" resultid="3976" />
                    <RANKING place="7" resultid="3979" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3" agemax="14" agemin="12" name="Jahrgang 2009 bis 2011">
                  <RANKINGS>
                    <RANKING place="7" resultid="26" />
                    <RANKING place="5" resultid="30" />
                    <RANKING place="11" resultid="576" />
                    <RANKING place="9" resultid="600" />
                    <RANKING place="1" resultid="1538" />
                    <RANKING place="10" resultid="1545" />
                    <RANKING place="17" resultid="1554" />
                    <RANKING place="12" resultid="1558" />
                    <RANKING place="8" resultid="1581" />
                    <RANKING place="6" resultid="2152" />
                    <RANKING place="3" resultid="2162" />
                    <RANKING place="4" resultid="2181" />
                    <RANKING place="14" resultid="3985" />
                    <RANKING place="16" resultid="4008" />
                    <RANKING place="15" resultid="4011" />
                    <RANKING place="13" resultid="4014" />
                    <RANKING place="2" resultid="4181" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="17" agemin="15" name="Jahrgang 2006 bis 2008">
                  <RANKINGS>
                    <RANKING place="8" resultid="584" />
                    <RANKING place="1" resultid="1560" />
                    <RANKING place="2" resultid="1578" />
                    <RANKING place="5" resultid="2171" />
                    <RANKING place="3" resultid="2175" />
                    <RANKING place="6" resultid="3988" />
                    <RANKING place="4" resultid="3998" />
                    <RANKING place="7" resultid="4002" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="42" number="104" gender="M" round="TIM">
              <SWIMSTYLE stroke="APNEA" name="25 Apnoe Männer" relaycount="1" distance="25" />
              <HEATS>
                <HEAT heatid="42001" number="1" />
                <HEAT heatid="42002" number="2" />
                <HEAT heatid="42003" number="3" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="2" agemax="11" agemin="10" name="Jahrgang 2012/2013">
                  <RANKINGS>
                    <RANKING place="5" resultid="570" />
                    <RANKING place="3" resultid="592" />
                    <RANKING place="7" resultid="607" />
                    <RANKING place="1" resultid="1541" />
                    <RANKING place="2" resultid="1550" />
                    <RANKING place="6" resultid="1592" />
                    <RANKING place="4" resultid="3982" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3" agemax="14" agemin="12" name="Jahrgang 2009 bis 2011">
                  <RANKINGS>
                    <RANKING place="1" resultid="2147" />
                    <RANKING place="3" resultid="2166" />
                    <RANKING place="2" resultid="2192" />
                    <RANKING place="4" resultid="4005" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="17" agemin="15" name="Jahrgang 2006 bis 2008">
                  <RANKINGS>
                    <RANKING place="4" resultid="1572" />
                    <RANKING place="2" resultid="1589" />
                    <RANKING place="3" resultid="1594" />
                    <RANKING place="1" resultid="2186" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="43" number="105" gender="F" round="TIM">
              <SWIMSTYLE stroke="SURFACE" name="25 Flossenschwimmen Frauen" relaycount="1" distance="25" />
              <HEATS>
                <HEAT heatid="43001" number="1" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="9" agemin="8" name="Jahrgang 2014/2015">
                  <RANKINGS>
                    <RANKING place="2" resultid="34" />
                    <RANKING place="3" resultid="42" />
                    <RANKING place="1" resultid="1586" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="44" number="106" gender="M" round="TIM">
              <SWIMSTYLE stroke="SURFACE" name="25 Flossenschwimmen Frauen" relaycount="1" distance="25" />
              <HEATS>
                <HEAT heatid="44001" number="1" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="9" agemin="8" name="Jahrgang 2014/2015">
                  <RANKINGS>
                    <RANKING place="3" resultid="38" />
                    <RANKING place="2" resultid="46" />
                    <RANKING place="1" resultid="588" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="7" number="7" gender="X" round="TIM">
              <SWIMSTYLE stroke="MEDLEY" relaycount="4" distance="50" />
              <HEATS>
                <HEAT heatid="7001" number="1" />
                <HEAT heatid="7002" number="2" />
                <HEAT heatid="7003" number="3" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="13" agemin="10" name="Jahrgang 2010 bis 2013">
                  <RANKINGS>
                    <RANKING place="2" resultid="111" />
                    <RANKING place="3" resultid="112" />
                    <RANKING place="5" resultid="3498" />
                    <RANKING place="19" resultid="3851" />
                    <RANKING place="13" resultid="4234" />
                    <RANKING place="11" resultid="4531" />
                    <RANKING place="8" resultid="4678" />
                    <RANKING place="14" resultid="4802" />
                    <RANKING place="18" resultid="4803" />
                    <RANKING place="6" resultid="5252" />
                    <RANKING place="7" resultid="5253" />
                    <RANKING place="15" resultid="5254" />
                    <RANKING place="4" resultid="5420" />
                    <RANKING place="12" resultid="5422" />
                    <RANKING place="1" resultid="5821" />
                    <RANKING place="9" resultid="5823" />
                    <RANKING place="10" resultid="5824" />
                    <RANKING place="16" resultid="5825" />
                    <RANKING place="17" resultid="5826" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
          </EVENTS>
        </SESSION>
        <SESSION number="2" date="2023-07-01" daytime="00:45">
          <EVENTS>
            <EVENT eventid="45" number="107" gender="F" round="TIM">
              <SWIMSTYLE stroke="SURFACE" name="100 Flossenschwimmen Frauen" relaycount="1" distance="100" />
              <HEATS>
                <HEAT heatid="45001" number="1" />
                <HEAT heatid="45002" number="2" />
                <HEAT heatid="45003" number="3" />
                <HEAT heatid="45004" number="4" />
                <HEAT heatid="45005" number="5" />
                <HEAT heatid="45006" number="6" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="9" agemin="8" name="Jahrgang 2014/2015">
                  <RANKINGS>
                    <RANKING place="3" resultid="35" />
                    <RANKING place="2" resultid="43" />
                    <RANKING place="1" resultid="1585" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2" agemax="11" agemin="10" name="Jahrgang 2012/2013">
                  <RANKINGS>
                    <RANKING place="5" resultid="581" />
                    <RANKING place="3" resultid="1530" />
                    <RANKING place="1" resultid="1562" />
                    <RANKING place="2" resultid="1566" />
                    <RANKING place="7" resultid="1575" />
                    <RANKING place="8" resultid="2168" />
                    <RANKING place="9" resultid="2178" />
                    <RANKING place="4" resultid="3977" />
                    <RANKING place="6" resultid="3980" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3" agemax="14" agemin="12" name="Jahrgang 2009 bis 2011">
                  <RANKINGS>
                    <RANKING place="6" resultid="27" />
                    <RANKING place="2" resultid="31" />
                    <RANKING place="18" resultid="574" />
                    <RANKING place="14" resultid="577" />
                    <RANKING place="8" resultid="601" />
                    <RANKING place="9" resultid="1544" />
                    <RANKING place="17" resultid="1553" />
                    <RANKING place="15" resultid="1557" />
                    <RANKING place="3" resultid="1580" />
                    <RANKING place="4" resultid="2151" />
                    <RANKING place="7" resultid="2161" />
                    <RANKING place="5" resultid="2180" />
                    <RANKING place="16" resultid="3971" />
                    <RANKING place="10" resultid="3986" />
                    <RANKING place="13" resultid="4009" />
                    <RANKING place="12" resultid="4012" />
                    <RANKING place="11" resultid="4015" />
                    <RANKING place="1" resultid="4182" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="17" agemin="15" name="Jahrgang 2006 bis 2008">
                  <RANKINGS>
                    <RANKING place="6" resultid="585" />
                    <RANKING place="10" resultid="597" />
                    <RANKING place="2" resultid="1534" />
                    <RANKING place="3" resultid="2170" />
                    <RANKING place="1" resultid="2174" />
                    <RANKING place="5" resultid="3989" />
                    <RANKING place="9" resultid="3992" />
                    <RANKING place="4" resultid="3999" />
                    <RANKING place="8" resultid="4003" />
                    <RANKING place="7" resultid="4018" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="46" number="108" gender="M" round="TIM">
              <SWIMSTYLE stroke="SURFACE" name="100 Flossenschwimmen Männer" relaycount="1" distance="100" />
              <HEATS>
                <HEAT heatid="46001" number="1" />
                <HEAT heatid="46002" number="2" />
                <HEAT heatid="46003" number="3" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="9" agemin="8" name="Jahrgang 2014/2015">
                  <RANKINGS>
                    <RANKING place="3" resultid="39" />
                    <RANKING place="2" resultid="47" />
                    <RANKING place="1" resultid="589" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2" agemax="11" agemin="10" name="Jahrgang 2012/2013">
                  <RANKINGS>
                    <RANKING place="8" resultid="567" />
                    <RANKING place="7" resultid="571" />
                    <RANKING place="4" resultid="593" />
                    <RANKING place="6" resultid="608" />
                    <RANKING place="1" resultid="1540" />
                    <RANKING place="3" resultid="1549" />
                    <RANKING place="5" resultid="2155" />
                    <RANKING place="9" resultid="2188" />
                    <RANKING place="2" resultid="3983" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3" agemax="14" agemin="12" name="Jahrgang 2009 bis 2011">
                  <RANKINGS>
                    <RANKING place="1" resultid="2146" />
                    <RANKING place="3" resultid="2158" />
                    <RANKING place="6" resultid="2165" />
                    <RANKING place="2" resultid="2191" />
                    <RANKING place="5" resultid="3974" />
                    <RANKING place="4" resultid="4006" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="17" agemin="15" name="Jahrgang 2006 bis 2008">
                  <RANKINGS>
                    <RANKING place="5" resultid="604" />
                    <RANKING place="4" resultid="1571" />
                    <RANKING place="1" resultid="1588" />
                    <RANKING place="3" resultid="1593" />
                    <RANKING place="2" resultid="2185" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="8" number="8" gender="F" round="TIM">
              <SWIMSTYLE stroke="FLY" relaycount="1" distance="200" />
              <HEATS>
                <HEAT heatid="8001" number="1" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="2" agemax="11" agemin="11" name="Jahrgang 2012">
                  <RANKINGS>
                    <RANKING place="1" resultid="5230" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="13" agemin="12" name="Jahrgang 2010/2011">
                  <RANKINGS>
                    <RANKING place="1" resultid="235" />
                    <RANKING place="2" resultid="2141" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6" agemax="15" agemin="14" name="Jahrgang 2008/2009">
                  <RANKINGS>
                    <RANKING place="1" resultid="5665" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8" agemax="17" agemin="16" name="Jahrgang 2006/2007">
                  <RANKINGS>
                    <RANKING place="1" resultid="5011" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="9" number="9" gender="M" round="TIM">
              <SWIMSTYLE stroke="FLY" relaycount="1" distance="200" />
              <HEATS>
                <HEAT heatid="9001" number="1" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="2" agemax="11" agemin="11" name="Jahrgang 2012" />
                <AGEGROUP agegroupid="4" agemax="13" agemin="12" name="Jahrgang 2010/2011">
                  <RANKINGS>
                    <RANKING place="2" resultid="241" />
                    <RANKING place="1" resultid="873" />
                    <RANKING place="4" resultid="1961" />
                    <RANKING place="3" resultid="6221" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6" agemax="15" agemin="14" name="Jahrgang 2008/2009" />
                <AGEGROUP agegroupid="8" agemax="17" agemin="16" name="Jahrgang 2006/2007" />
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="10" number="10" gender="F" round="TIM">
              <SWIMSTYLE stroke="BACK" relaycount="1" distance="100" />
              <HEATS>
                <HEAT heatid="10001" number="1" />
                <HEAT heatid="10002" number="2" />
                <HEAT heatid="10003" number="3" />
                <HEAT heatid="10004" number="4" />
                <HEAT heatid="10005" number="5" />
                <HEAT heatid="10006" number="6" />
                <HEAT heatid="10007" number="7" />
                <HEAT heatid="10008" number="8" />
                <HEAT heatid="10009" number="9" />
                <HEAT heatid="10010" number="10" />
                <HEAT heatid="10011" number="11" />
                <HEAT heatid="10012" number="12" />
                <HEAT heatid="10013" number="13" />
                <HEAT heatid="10014" number="14" />
                <HEAT heatid="10015" number="15" />
                <HEAT heatid="10016" number="16" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="10" agemin="10" name="Jahrgang 2013">
                  <RANKINGS>
                    <RANKING place="3" resultid="9" />
                    <RANKING place="9" resultid="208" />
                    <RANKING place="6" resultid="242" />
                    <RANKING place="11" resultid="844" />
                    <RANKING place="5" resultid="890" />
                    <RANKING place="16" resultid="952" />
                    <RANKING place="7" resultid="1921" />
                    <RANKING place="10" resultid="2122" />
                    <RANKING place="18" resultid="3731" />
                    <RANKING place="20" resultid="4126" />
                    <RANKING place="15" resultid="4158" />
                    <RANKING place="19" resultid="4261" />
                    <RANKING place="14" resultid="4633" />
                    <RANKING place="17" resultid="4958" />
                    <RANKING place="1" resultid="5140" />
                    <RANKING place="12" resultid="5190" />
                    <RANKING place="8" resultid="5219" />
                    <RANKING place="4" resultid="5440" />
                    <RANKING place="2" resultid="5574" />
                    <RANKING place="13" resultid="6048" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2" agemax="11" agemin="11" name="Jahrgang 2012">
                  <RANKINGS>
                    <RANKING place="11" resultid="16" />
                    <RANKING place="14" resultid="179" />
                    <RANKING place="12" resultid="959" />
                    <RANKING place="17" resultid="1610" />
                    <RANKING place="19" resultid="1616" />
                    <RANKING place="29" resultid="1653" />
                    <RANKING place="9" resultid="1994" />
                    <RANKING place="22" resultid="2115" />
                    <RANKING place="8" resultid="2125" />
                    <RANKING place="31" resultid="4320" />
                    <RANKING place="13" resultid="4501" />
                    <RANKING place="4" resultid="4505" />
                    <RANKING place="5" resultid="4738" />
                    <RANKING place="21" resultid="4811" />
                    <RANKING place="34" resultid="4872" />
                    <RANKING place="10" resultid="4911" />
                    <RANKING place="23" resultid="4918" />
                    <RANKING place="33" resultid="5106" />
                    <RANKING place="27" resultid="5178" />
                    <RANKING place="2" resultid="5342" />
                    <RANKING place="25" resultid="5491" />
                    <RANKING place="36" resultid="5616" />
                    <RANKING place="15" resultid="5643" />
                    <RANKING place="32" resultid="5670" />
                    <RANKING place="3" resultid="5711" />
                    <RANKING place="24" resultid="5719" />
                    <RANKING place="35" resultid="5794" />
                    <RANKING place="6" resultid="5842" />
                    <RANKING place="18" resultid="5931" />
                    <RANKING place="26" resultid="5973" />
                    <RANKING place="7" resultid="6035" />
                    <RANKING place="1" resultid="6064" />
                    <RANKING place="28" resultid="6177" />
                    <RANKING place="20" resultid="6317" />
                    <RANKING place="30" resultid="6337" />
                    <RANKING place="16" resultid="6345" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="13" agemin="12" name="Jahrgang 2010/2011">
                  <RANKINGS>
                    <RANKING place="23" resultid="147" />
                    <RANKING place="9" resultid="155" />
                    <RANKING place="10" resultid="171" />
                    <RANKING place="11" resultid="218" />
                    <RANKING place="4" resultid="613" />
                    <RANKING place="6" resultid="976" />
                    <RANKING place="20" resultid="1947" />
                    <RANKING place="21" resultid="2063" />
                    <RANKING place="1" resultid="3453" />
                    <RANKING place="32" resultid="3742" />
                    <RANKING place="25" resultid="3762" />
                    <RANKING place="33" resultid="3781" />
                    <RANKING place="12" resultid="4061" />
                    <RANKING place="31" resultid="4108" />
                    <RANKING place="15" resultid="4388" />
                    <RANKING place="7" resultid="4440" />
                    <RANKING place="29" resultid="4557" />
                    <RANKING place="18" resultid="4865" />
                    <RANKING place="28" resultid="4878" />
                    <RANKING place="14" resultid="4928" />
                    <RANKING place="21" resultid="5084" />
                    <RANKING place="19" resultid="5146" />
                    <RANKING place="8" resultid="5207" />
                    <RANKING place="5" resultid="5238" />
                    <RANKING place="27" resultid="5280" />
                    <RANKING place="13" resultid="5328" />
                    <RANKING place="3" resultid="5391" />
                    <RANKING place="16" resultid="5403" />
                    <RANKING place="26" resultid="5759" />
                    <RANKING place="17" resultid="5788" />
                    <RANKING place="30" resultid="6078" />
                    <RANKING place="2" resultid="6114" />
                    <RANKING place="24" resultid="6283" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6" agemax="15" agemin="14" name="Jahrgang 2008/2009">
                  <RANKINGS>
                    <RANKING place="1" resultid="2012" />
                    <RANKING place="13" resultid="3463" />
                    <RANKING place="7" resultid="3473" />
                    <RANKING place="2" resultid="4579" />
                    <RANKING place="6" resultid="4941" />
                    <RANKING place="3" resultid="4994" />
                    <RANKING place="11" resultid="5059" />
                    <RANKING place="12" resultid="5321" />
                    <RANKING place="4" resultid="5353" />
                    <RANKING place="14" resultid="5455" />
                    <RANKING place="10" resultid="5733" />
                    <RANKING place="8" resultid="5919" />
                    <RANKING place="9" resultid="6157" />
                    <RANKING place="5" resultid="6275" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8" agemax="17" agemin="16" name="Jahrgang 2006/2007">
                  <RANKINGS>
                    <RANKING place="8" resultid="1911" />
                    <RANKING place="7" resultid="4622" />
                    <RANKING place="6" resultid="4649" />
                    <RANKING place="1" resultid="4673" />
                    <RANKING place="3" resultid="4702" />
                    <RANKING place="5" resultid="5012" />
                    <RANKING place="2" resultid="5487" />
                    <RANKING place="4" resultid="6351" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="11" number="11" gender="M" round="TIM">
              <SWIMSTYLE stroke="BACK" relaycount="1" distance="100" />
              <HEATS>
                <HEAT heatid="11001" number="1" />
                <HEAT heatid="11002" number="2" />
                <HEAT heatid="11003" number="3" />
                <HEAT heatid="11004" number="4" />
                <HEAT heatid="11005" number="5" />
                <HEAT heatid="11006" number="6" />
                <HEAT heatid="11007" number="7" />
                <HEAT heatid="11008" number="8" />
                <HEAT heatid="11009" number="9" />
                <HEAT heatid="11010" number="10" />
                <HEAT heatid="11011" number="11" />
                <HEAT heatid="11012" number="12" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="10" agemin="10" name="Jahrgang 2013">
                  <RANKINGS>
                    <RANKING place="1" resultid="945" />
                    <RANKING place="10" resultid="1626" />
                    <RANKING place="3" resultid="3438" />
                    <RANKING place="15" resultid="3806" />
                    <RANKING place="12" resultid="4175" />
                    <RANKING place="13" resultid="4247" />
                    <RANKING place="8" resultid="4758" />
                    <RANKING place="9" resultid="4776" />
                    <RANKING place="2" resultid="4982" />
                    <RANKING place="14" resultid="5062" />
                    <RANKING place="4" resultid="5260" />
                    <RANKING place="11" resultid="5585" />
                    <RANKING place="6" resultid="5887" />
                    <RANKING place="7" resultid="6197" />
                    <RANKING place="5" resultid="6260" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2" agemax="11" agemin="11" name="Jahrgang 2012">
                  <RANKINGS>
                    <RANKING place="2" resultid="123" />
                    <RANKING place="1" resultid="187" />
                    <RANKING place="7" resultid="822" />
                    <RANKING place="23" resultid="859" />
                    <RANKING place="17" resultid="917" />
                    <RANKING place="20" resultid="993" />
                    <RANKING place="27" resultid="1001" />
                    <RANKING place="10" resultid="2009" />
                    <RANKING place="4" resultid="2107" />
                    <RANKING place="28" resultid="2111" />
                    <RANKING place="13" resultid="2118" />
                    <RANKING place="24" resultid="4065" />
                    <RANKING place="11" resultid="4111" />
                    <RANKING place="29" resultid="4168" />
                    <RANKING place="18" resultid="4267" />
                    <RANKING place="21" resultid="4717" />
                    <RANKING place="5" resultid="4724" />
                    <RANKING place="15" resultid="4796" />
                    <RANKING place="3" resultid="5169" />
                    <RANKING place="22" resultid="5306" />
                    <RANKING place="6" resultid="5517" />
                    <RANKING place="8" resultid="5524" />
                    <RANKING place="25" resultid="5566" />
                    <RANKING place="9" resultid="5686" />
                    <RANKING place="16" resultid="5802" />
                    <RANKING place="19" resultid="5849" />
                    <RANKING place="12" resultid="5939" />
                    <RANKING place="26" resultid="6100" />
                    <RANKING place="14" resultid="6293" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="13" agemin="12" name="Jahrgang 2010/2011">
                  <RANKINGS>
                    <RANKING place="2" resultid="115" />
                    <RANKING place="6" resultid="139" />
                    <RANKING place="3" resultid="794" />
                    <RANKING place="10" resultid="1933" />
                    <RANKING place="9" resultid="1938" />
                    <RANKING place="19" resultid="2024" />
                    <RANKING place="14" resultid="2092" />
                    <RANKING place="18" resultid="3476" />
                    <RANKING place="4" resultid="4022" />
                    <RANKING place="12" resultid="4076" />
                    <RANKING place="1" resultid="4466" />
                    <RANKING place="17" resultid="4540" />
                    <RANKING place="25" resultid="4569" />
                    <RANKING place="15" resultid="4591" />
                    <RANKING place="20" resultid="4604" />
                    <RANKING place="24" resultid="4609" />
                    <RANKING place="22" resultid="4639" />
                    <RANKING place="7" resultid="4791" />
                    <RANKING place="21" resultid="4898" />
                    <RANKING place="23" resultid="5264" />
                    <RANKING place="16" resultid="5284" />
                    <RANKING place="8" resultid="5424" />
                    <RANKING place="5" resultid="5747" />
                    <RANKING place="11" resultid="5881" />
                    <RANKING place="26" resultid="6031" />
                    <RANKING place="13" resultid="6328" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6" agemax="15" agemin="14" name="Jahrgang 2008/2009">
                  <RANKINGS>
                    <RANKING place="7" resultid="231" />
                    <RANKING place="5" resultid="3835" />
                    <RANKING place="3" resultid="4597" />
                    <RANKING place="6" resultid="4819" />
                    <RANKING place="2" resultid="4851" />
                    <RANKING place="4" resultid="4905" />
                    <RANKING place="1" resultid="5386" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8" agemax="17" agemin="16" name="Jahrgang 2006/2007">
                  <RANKINGS>
                    <RANKING place="2" resultid="3467" />
                    <RANKING place="6" resultid="3486" />
                    <RANKING place="5" resultid="4575" />
                    <RANKING place="3" resultid="4708" />
                    <RANKING place="4" resultid="5133" />
                    <RANKING place="1" resultid="5314" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="47" number="109" gender="F" round="TIM">
              <SWIMSTYLE stroke="UNKNOWN" name="50 Torstoß Frauen" relaycount="1" distance="50" />
              <HEATS>
                <HEAT heatid="47001" number="1" />
                <HEAT heatid="47002" number="2" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="11" agemin="8" name="Kategorie U12">
                  <RANKINGS>
                    <RANKING place="3" resultid="1529" />
                    <RANKING place="1" resultid="1561" />
                    <RANKING place="4" resultid="1565" />
                    <RANKING place="2" resultid="1574" />
                    <RANKING place="5" resultid="1584" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2" agemax="14" agemin="12" name="Kategorie U15">
                  <RANKINGS>
                    <RANKING place="1" resultid="1537" />
                    <RANKING place="4" resultid="1543" />
                    <RANKING place="5" resultid="1552" />
                    <RANKING place="6" resultid="1556" />
                    <RANKING place="2" resultid="1579" />
                    <RANKING place="3" resultid="2150" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3" agemax="17" agemin="15" name="Kategorie U18">
                  <RANKINGS>
                    <RANKING place="1" resultid="1533" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="48" number="110" gender="M" round="TIM">
              <SWIMSTYLE stroke="UNKNOWN" name="50 Torstoß Männer" relaycount="1" distance="50" />
              <HEATS>
                <HEAT heatid="48001" number="1" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="11" agemin="8" name="Kategorie U12">
                  <RANKINGS>
                    <RANKING place="1" resultid="1539" />
                    <RANKING place="2" resultid="1548" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2" agemax="14" agemin="12" name="Kategorie U15">
                  <RANKINGS>
                    <RANKING place="2" resultid="2145" />
                    <RANKING place="1" resultid="2164" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3" agemax="17" agemin="15" name="Kategorie U18">
                  <RANKINGS>
                    <RANKING place="3" resultid="1570" />
                    <RANKING place="2" resultid="1587" />
                    <RANKING place="1" resultid="2184" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="12" number="12" gender="F" round="TIM">
              <SWIMSTYLE stroke="FREE" relaycount="1" distance="50" />
              <HEATS>
                <HEAT heatid="12001" number="1" />
                <HEAT heatid="12002" number="2" />
                <HEAT heatid="12003" number="3" />
                <HEAT heatid="12004" number="4" />
                <HEAT heatid="12005" number="5" />
                <HEAT heatid="12006" number="6" />
                <HEAT heatid="12007" number="7" />
                <HEAT heatid="12008" number="8" />
                <HEAT heatid="12009" number="9" />
                <HEAT heatid="12010" number="10" />
                <HEAT heatid="12011" number="11" />
                <HEAT heatid="12012" number="12" />
                <HEAT heatid="12013" number="13" />
                <HEAT heatid="12014" number="14" />
                <HEAT heatid="12015" number="15" />
                <HEAT heatid="12016" number="16" />
                <HEAT heatid="12017" number="17" />
                <HEAT heatid="12018" number="18" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="10" agemin="10" name="Jahrgang 2013">
                  <RANKINGS>
                    <RANKING place="4" resultid="10" />
                    <RANKING place="2" resultid="209" />
                    <RANKING place="8" resultid="243" />
                    <RANKING place="6" resultid="472" />
                    <RANKING place="10" resultid="843" />
                    <RANKING place="5" resultid="889" />
                    <RANKING place="11" resultid="897" />
                    <RANKING place="28" resultid="951" />
                    <RANKING place="13" resultid="1920" />
                    <RANKING place="7" resultid="2121" />
                    <RANKING place="19" resultid="3730" />
                    <RANKING place="23" resultid="4127" />
                    <RANKING place="26" resultid="4159" />
                    <RANKING place="27" resultid="4257" />
                    <RANKING place="22" resultid="4262" />
                    <RANKING place="12" resultid="4616" />
                    <RANKING place="20" resultid="4634" />
                    <RANKING place="16" resultid="4690" />
                    <RANKING place="14" resultid="4747" />
                    <RANKING place="18" resultid="4959" />
                    <RANKING place="25" resultid="5095" />
                    <RANKING place="2" resultid="5141" />
                    <RANKING place="24" resultid="5162" />
                    <RANKING place="15" resultid="5191" />
                    <RANKING place="1" resultid="5441" />
                    <RANKING place="9" resultid="5575" />
                    <RANKING place="17" resultid="5829" />
                    <RANKING place="21" resultid="6049" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2" agemax="11" agemin="11" name="Jahrgang 2012">
                  <RANKINGS>
                    <RANKING place="3" resultid="17" />
                    <RANKING place="13" resultid="180" />
                    <RANKING place="5" resultid="958" />
                    <RANKING place="16" resultid="1598" />
                    <RANKING place="17" resultid="1609" />
                    <RANKING place="12" resultid="1615" />
                    <RANKING place="33" resultid="1647" />
                    <RANKING place="28" resultid="1652" />
                    <RANKING place="14" resultid="1895" />
                    <RANKING place="27" resultid="1953" />
                    <RANKING place="7" resultid="1993" />
                    <RANKING place="25" resultid="2114" />
                    <RANKING place="10" resultid="2124" />
                    <RANKING place="20" resultid="4321" />
                    <RANKING place="2" resultid="4436" />
                    <RANKING place="8" resultid="4739" />
                    <RANKING place="19" resultid="4812" />
                    <RANKING place="23" resultid="4858" />
                    <RANKING place="29" resultid="4873" />
                    <RANKING place="18" resultid="4912" />
                    <RANKING place="24" resultid="4919" />
                    <RANKING place="26" resultid="5035" />
                    <RANKING place="35" resultid="5107" />
                    <RANKING place="9" resultid="5179" />
                    <RANKING place="15" resultid="5231" />
                    <RANKING place="34" resultid="5617" />
                    <RANKING place="4" resultid="5712" />
                    <RANKING place="31" resultid="5795" />
                    <RANKING place="22" resultid="5843" />
                    <RANKING place="21" resultid="5932" />
                    <RANKING place="32" resultid="6023" />
                    <RANKING place="11" resultid="6036" />
                    <RANKING place="1" resultid="6065" />
                    <RANKING place="30" resultid="6338" />
                    <RANKING place="6" resultid="6364" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="13" agemin="12" name="Jahrgang 2010/2011">
                  <RANKINGS>
                    <RANKING place="4" resultid="131" />
                    <RANKING place="8" resultid="156" />
                    <RANKING place="5" resultid="172" />
                    <RANKING place="3" resultid="614" />
                    <RANKING place="14" resultid="975" />
                    <RANKING place="19" resultid="1946" />
                    <RANKING place="15" resultid="1989" />
                    <RANKING place="24" resultid="2062" />
                    <RANKING place="9" resultid="2140" />
                    <RANKING place="39" resultid="3741" />
                    <RANKING place="17" resultid="4030" />
                    <RANKING place="6" resultid="4062" />
                    <RANKING place="33" resultid="4109" />
                    <RANKING place="31" resultid="4133" />
                    <RANKING place="21" resultid="4389" />
                    <RANKING place="12" resultid="4441" />
                    <RANKING place="26" resultid="4546" />
                    <RANKING place="38" resultid="4558" />
                    <RANKING place="13" resultid="4866" />
                    <RANKING place="25" resultid="4879" />
                    <RANKING place="20" resultid="4929" />
                    <RANKING place="36" resultid="5001" />
                    <RANKING place="23" resultid="5085" />
                    <RANKING place="27" resultid="5147" />
                    <RANKING place="16" resultid="5208" />
                    <RANKING place="10" resultid="5239" />
                    <RANKING place="7" resultid="5256" />
                    <RANKING place="35" resultid="5281" />
                    <RANKING place="22" resultid="5462" />
                    <RANKING place="1" resultid="5500" />
                    <RANKING place="30" resultid="5606" />
                    <RANKING place="37" resultid="5706" />
                    <RANKING place="34" resultid="5760" />
                    <RANKING place="32" resultid="5775" />
                    <RANKING place="29" resultid="5786" />
                    <RANKING place="18" resultid="5789" />
                    <RANKING place="11" resultid="5800" />
                    <RANKING place="41" resultid="6004" />
                    <RANKING place="40" resultid="6079" />
                    <RANKING place="2" resultid="6137" />
                    <RANKING place="28" resultid="6284" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6" agemax="15" agemin="14" name="Jahrgang 2008/2009">
                  <RANKINGS>
                    <RANKING place="19" resultid="3462" />
                    <RANKING place="12" resultid="3472" />
                    <RANKING place="10" resultid="3722" />
                    <RANKING place="4" resultid="4580" />
                    <RANKING place="17" resultid="4743" />
                    <RANKING place="13" resultid="4886" />
                    <RANKING place="5" resultid="4942" />
                    <RANKING place="7" resultid="4995" />
                    <RANKING place="8" resultid="5060" />
                    <RANKING place="2" resultid="5354" />
                    <RANKING place="3" resultid="5432" />
                    <RANKING place="16" resultid="5456" />
                    <RANKING place="9" resultid="5609" />
                    <RANKING place="15" resultid="5734" />
                    <RANKING place="14" resultid="5874" />
                    <RANKING place="11" resultid="5914" />
                    <RANKING place="18" resultid="5920" />
                    <RANKING place="1" resultid="6042" />
                    <RANKING place="6" resultid="6276" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8" agemax="17" agemin="16" name="Jahrgang 2006/2007">
                  <RANKINGS>
                    <RANKING place="6" resultid="1910" />
                    <RANKING place="3" resultid="4623" />
                    <RANKING place="4" resultid="4650" />
                    <RANKING place="5" resultid="4730" />
                    <RANKING place="7" resultid="4839" />
                    <RANKING place="8" resultid="5013" />
                    <RANKING place="1" resultid="6161" />
                    <RANKING place="2" resultid="6352" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="13" number="13" gender="M" round="TIM">
              <SWIMSTYLE stroke="FREE" relaycount="1" distance="50" />
              <HEATS>
                <HEAT heatid="13001" number="1" />
                <HEAT heatid="13002" number="2" />
                <HEAT heatid="13003" number="3" />
                <HEAT heatid="13004" number="4" />
                <HEAT heatid="13005" number="5" />
                <HEAT heatid="13006" number="6" />
                <HEAT heatid="13007" number="7" />
                <HEAT heatid="13008" number="8" />
                <HEAT heatid="13009" number="9" />
                <HEAT heatid="13010" number="10" />
                <HEAT heatid="13011" number="11" />
                <HEAT heatid="13012" number="12" />
                <HEAT heatid="13013" number="13" />
                <HEAT heatid="13014" number="14" />
                <HEAT heatid="13015" number="15" />
                <HEAT heatid="13016" number="16" />
                <HEAT heatid="13017" number="17" />
                <HEAT heatid="13018" number="18" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="10" agemin="10" name="Jahrgang 2013">
                  <RANKINGS>
                    <RANKING place="8" resultid="829" />
                    <RANKING place="6" resultid="852" />
                    <RANKING place="3" resultid="944" />
                    <RANKING place="16" resultid="1632" />
                    <RANKING place="1" resultid="3437" />
                    <RANKING place="24" resultid="3803" />
                    <RANKING place="25" resultid="3805" />
                    <RANKING place="5" resultid="4039" />
                    <RANKING place="7" resultid="4051" />
                    <RANKING place="12" resultid="4098" />
                    <RANKING place="11" resultid="4176" />
                    <RANKING place="14" resultid="4248" />
                    <RANKING place="9" resultid="4759" />
                    <RANKING place="15" resultid="4777" />
                    <RANKING place="13" resultid="4983" />
                    <RANKING place="21" resultid="5063" />
                    <RANKING place="18" resultid="5261" />
                    <RANKING place="23" resultid="5337" />
                    <RANKING place="10" resultid="5586" />
                    <RANKING place="2" resultid="5625" />
                    <RANKING place="20" resultid="5888" />
                    <RANKING place="4" resultid="5951" />
                    <RANKING place="22" resultid="6127" />
                    <RANKING place="19" resultid="6198" />
                    <RANKING place="17" resultid="6261" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2" agemax="11" agemin="11" name="Jahrgang 2012">
                  <RANKINGS>
                    <RANKING place="2" resultid="124" />
                    <RANKING place="25" resultid="163" />
                    <RANKING place="3" resultid="188" />
                    <RANKING place="22" resultid="814" />
                    <RANKING place="26" resultid="858" />
                    <RANKING place="11" resultid="916" />
                    <RANKING place="19" resultid="992" />
                    <RANKING place="27" resultid="1000" />
                    <RANKING place="7" resultid="2106" />
                    <RANKING place="28" resultid="2110" />
                    <RANKING place="17" resultid="2117" />
                    <RANKING place="33" resultid="3750" />
                    <RANKING place="32" resultid="3790" />
                    <RANKING place="12" resultid="4066" />
                    <RANKING place="8" resultid="4112" />
                    <RANKING place="31" resultid="4169" />
                    <RANKING place="14" resultid="4268" />
                    <RANKING place="20" resultid="4718" />
                    <RANKING place="6" resultid="4725" />
                    <RANKING place="16" resultid="4826" />
                    <RANKING place="10" resultid="5170" />
                    <RANKING place="21" resultid="5307" />
                    <RANKING place="9" resultid="5414" />
                    <RANKING place="5" resultid="5518" />
                    <RANKING place="15" resultid="5525" />
                    <RANKING place="34" resultid="5547" />
                    <RANKING place="23" resultid="5567" />
                    <RANKING place="4" resultid="5687" />
                    <RANKING place="24" resultid="5803" />
                    <RANKING place="35" resultid="5808" />
                    <RANKING place="29" resultid="5850" />
                    <RANKING place="18" resultid="5940" />
                    <RANKING place="30" resultid="6101" />
                    <RANKING place="1" resultid="6184" />
                    <RANKING place="13" resultid="6294" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="13" agemin="12" name="Jahrgang 2010/2011">
                  <RANKINGS>
                    <RANKING place="12" resultid="116" />
                    <RANKING place="10" resultid="140" />
                    <RANKING place="3" resultid="772" />
                    <RANKING place="7" resultid="793" />
                    <RANKING place="1" resultid="872" />
                    <RANKING place="25" resultid="1932" />
                    <RANKING place="18" resultid="1937" />
                    <RANKING place="33" resultid="2023" />
                    <RANKING place="35" resultid="2091" />
                    <RANKING place="15" resultid="3444" />
                    <RANKING place="23" resultid="3475" />
                    <RANKING place="38" resultid="3814" />
                    <RANKING place="40" resultid="3849" />
                    <RANKING place="9" resultid="4023" />
                    <RANKING place="30" resultid="4077" />
                    <RANKING place="14" resultid="4285" />
                    <RANKING place="8" resultid="4467" />
                    <RANKING place="29" resultid="4541" />
                    <RANKING place="22" resultid="4552" />
                    <RANKING place="36" resultid="4570" />
                    <RANKING place="6" resultid="4592" />
                    <RANKING place="19" resultid="4605" />
                    <RANKING place="31" resultid="4610" />
                    <RANKING place="2" resultid="4627" />
                    <RANKING place="37" resultid="4640" />
                    <RANKING place="5" resultid="4792" />
                    <RANKING place="20" resultid="4892" />
                    <RANKING place="34" resultid="4899" />
                    <RANKING place="27" resultid="5265" />
                    <RANKING place="32" resultid="5285" />
                    <RANKING place="17" resultid="5425" />
                    <RANKING place="16" resultid="5660" />
                    <RANKING place="4" resultid="5698" />
                    <RANKING place="28" resultid="5740" />
                    <RANKING place="11" resultid="5743" />
                    <RANKING place="13" resultid="5748" />
                    <RANKING place="26" resultid="5882" />
                    <RANKING place="23" resultid="5897" />
                    <RANKING place="39" resultid="6032" />
                    <RANKING place="41" resultid="6210" />
                    <RANKING place="21" resultid="6329" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6" agemax="15" agemin="14" name="Jahrgang 2008/2009">
                  <RANKINGS>
                    <RANKING place="19" resultid="3770" />
                    <RANKING place="3" resultid="4105" />
                    <RANKING place="2" resultid="4316" />
                    <RANKING place="20" resultid="4537" />
                    <RANKING place="16" resultid="4598" />
                    <RANKING place="11" resultid="4661" />
                    <RANKING place="8" resultid="4783" />
                    <RANKING place="15" resultid="4805" />
                    <RANKING place="17" resultid="4820" />
                    <RANKING place="10" resultid="4852" />
                    <RANKING place="7" resultid="4906" />
                    <RANKING place="8" resultid="4951" />
                    <RANKING place="18" resultid="5682" />
                    <RANKING place="13" resultid="5766" />
                    <RANKING place="4" resultid="5901" />
                    <RANKING place="6" resultid="5999" />
                    <RANKING place="1" resultid="6018" />
                    <RANKING place="12" resultid="6081" />
                    <RANKING place="14" resultid="6096" />
                    <RANKING place="5" resultid="6141" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8" agemax="17" agemin="16" name="Jahrgang 2006/2007">
                  <RANKINGS>
                    <RANKING place="3" resultid="3466" />
                    <RANKING place="7" resultid="3485" />
                    <RANKING place="10" resultid="3798" />
                    <RANKING place="11" resultid="4295" />
                    <RANKING place="5" resultid="4576" />
                    <RANKING place="1" resultid="4709" />
                    <RANKING place="9" resultid="4833" />
                    <RANKING place="4" resultid="5134" />
                    <RANKING place="2" resultid="5315" />
                    <RANKING place="8" resultid="5563" />
                    <RANKING place="6" resultid="5581" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="14" number="14" gender="F" round="TIM">
              <SWIMSTYLE stroke="BREAST" relaycount="1" distance="200" />
              <HEATS>
                <HEAT heatid="14001" number="1" />
                <HEAT heatid="14002" number="2" />
                <HEAT heatid="14003" number="3" />
                <HEAT heatid="14004" number="4" />
                <HEAT heatid="14005" number="5" />
                <HEAT heatid="14006" number="6" />
                <HEAT heatid="14007" number="7" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="10" agemin="10" name="Jahrgang 2013">
                  <RANKINGS>
                    <RANKING place="4" resultid="210" />
                    <RANKING place="5" resultid="244" />
                    <RANKING place="3" resultid="896" />
                    <RANKING place="7" resultid="3827" />
                    <RANKING place="10" resultid="4258" />
                    <RANKING place="8" resultid="4691" />
                    <RANKING place="6" resultid="4748" />
                    <RANKING place="1" resultid="5220" />
                    <RANKING place="9" resultid="5779" />
                    <RANKING place="2" resultid="5830" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2" agemax="11" agemin="11" name="Jahrgang 2012">
                  <RANKINGS>
                    <RANKING place="2" resultid="1894" />
                    <RANKING place="6" resultid="1952" />
                    <RANKING place="7" resultid="1956" />
                    <RANKING place="1" resultid="4437" />
                    <RANKING place="10" resultid="4502" />
                    <RANKING place="8" resultid="4506" />
                    <RANKING place="12" resultid="5492" />
                    <RANKING place="14" resultid="5618" />
                    <RANKING place="5" resultid="5644" />
                    <RANKING place="13" resultid="5671" />
                    <RANKING place="11" resultid="5720" />
                    <RANKING place="9" resultid="6024" />
                    <RANKING place="4" resultid="6318" />
                    <RANKING place="3" resultid="6346" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="13" agemin="12" name="Jahrgang 2010/2011">
                  <RANKINGS>
                    <RANKING place="1" resultid="132" />
                    <RANKING place="4" resultid="148" />
                    <RANKING place="11" resultid="1988" />
                    <RANKING place="5" resultid="3761" />
                    <RANKING place="8" resultid="4031" />
                    <RANKING place="16" resultid="4110" />
                    <RANKING place="12" resultid="4547" />
                    <RANKING place="15" resultid="4696" />
                    <RANKING place="6" resultid="4880" />
                    <RANKING place="7" resultid="5257" />
                    <RANKING place="9" resultid="5369" />
                    <RANKING place="3" resultid="5392" />
                    <RANKING place="2" resultid="5437" />
                    <RANKING place="18" resultid="5503" />
                    <RANKING place="17" resultid="5761" />
                    <RANKING place="10" resultid="5776" />
                    <RANKING place="14" resultid="6005" />
                    <RANKING place="13" resultid="6361" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6" agemax="15" agemin="14" name="Jahrgang 2008/2009">
                  <RANKINGS>
                    <RANKING place="3" resultid="3822" />
                    <RANKING place="2" resultid="5497" />
                    <RANKING place="4" resultid="5650" />
                    <RANKING place="1" resultid="5877" />
                    <RANKING place="5" resultid="6189" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8" agemax="17" agemin="16" name="Jahrgang 2006/2007">
                  <RANKINGS>
                    <RANKING place="2" resultid="4624" />
                    <RANKING place="1" resultid="4703" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="15" number="15" gender="M" round="TIM">
              <SWIMSTYLE stroke="BREAST" relaycount="1" distance="200" />
              <HEATS>
                <HEAT heatid="15001" number="1" />
                <HEAT heatid="15002" number="2" />
                <HEAT heatid="15003" number="3" />
                <HEAT heatid="15004" number="4" />
                <HEAT heatid="15005" number="5" />
                <HEAT heatid="15006" number="6" />
                <HEAT heatid="15007" number="7" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="10" agemin="10" name="Jahrgang 2013">
                  <RANKINGS>
                    <RANKING place="4" resultid="851" />
                    <RANKING place="7" resultid="1625" />
                    <RANKING place="1" resultid="1631" />
                    <RANKING place="2" resultid="4040" />
                    <RANKING place="8" resultid="4099" />
                    <RANKING place="6" resultid="4760" />
                    <RANKING place="9" resultid="5338" />
                    <RANKING place="3" resultid="5587" />
                    <RANKING place="5" resultid="5952" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2" agemax="11" agemin="11" name="Jahrgang 2012">
                  <RANKINGS>
                    <RANKING place="10" resultid="164" />
                    <RANKING place="4" resultid="821" />
                    <RANKING place="5" resultid="2008" />
                    <RANKING place="1" resultid="3458" />
                    <RANKING place="2" resultid="4113" />
                    <RANKING place="7" resultid="4797" />
                    <RANKING place="6" resultid="5308" />
                    <RANKING place="8" resultid="5526" />
                    <RANKING place="11" resultid="5548" />
                    <RANKING place="12" resultid="5809" />
                    <RANKING place="3" resultid="5816" />
                    <RANKING place="9" resultid="6102" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="13" agemin="12" name="Jahrgang 2010/2011">
                  <RANKINGS>
                    <RANKING place="2" resultid="771" />
                    <RANKING place="3" resultid="3443" />
                    <RANKING place="10" resultid="3813" />
                    <RANKING place="8" resultid="4078" />
                    <RANKING place="4" resultid="4628" />
                    <RANKING place="5" resultid="4793" />
                    <RANKING place="11" resultid="4900" />
                    <RANKING place="7" resultid="5273" />
                    <RANKING place="1" resultid="5453" />
                    <RANKING place="9" resultid="5741" />
                    <RANKING place="6" resultid="5744" />
                    <RANKING place="12" resultid="6211" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6" agemax="15" agemin="14" name="Jahrgang 2008/2009">
                  <RANKINGS>
                    <RANKING place="10" resultid="233" />
                    <RANKING place="6" resultid="3715" />
                    <RANKING place="3" resultid="3776" />
                    <RANKING place="9" resultid="4106" />
                    <RANKING place="8" resultid="4599" />
                    <RANKING place="2" resultid="4784" />
                    <RANKING place="11" resultid="4806" />
                    <RANKING place="5" resultid="4952" />
                    <RANKING place="4" resultid="5361" />
                    <RANKING place="7" resultid="5767" />
                    <RANKING place="1" resultid="5836" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8" agemax="17" agemin="16" name="Jahrgang 2006/2007">
                  <RANKINGS>
                    <RANKING place="1" resultid="4296" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="16" number="16" gender="X" round="TIM">
              <SWIMSTYLE stroke="MEDLEY" relaycount="4" distance="50" />
              <HEATS>
                <HEAT heatid="16001" number="1" />
                <HEAT heatid="16002" number="2" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="17" agemin="14" name="Jahrgang 2006 bis 2009">
                  <RANKINGS>
                    <RANKING place="4" resultid="3499" />
                    <RANKING place="7" resultid="4530" />
                    <RANKING place="5" resultid="4677" />
                    <RANKING place="6" resultid="4801" />
                    <RANKING place="3" resultid="5251" />
                    <RANKING place="2" resultid="5419" />
                    <RANKING place="8" resultid="5421" />
                    <RANKING place="1" resultid="5822" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="49" number="111" gender="F" round="TIM">
              <SWIMSTYLE stroke="SURFACE" name="50 Flossenschwimmen Frauen" relaycount="1" distance="50" />
              <HEATS>
                <HEAT heatid="49001" number="1" />
                <HEAT heatid="49002" number="2" />
                <HEAT heatid="49003" number="3" />
                <HEAT heatid="49004" number="4" />
                <HEAT heatid="49005" number="5" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="9" agemin="8" name="Jahrgang 2014/2015">
                  <RANKINGS>
                    <RANKING place="3" resultid="36" />
                    <RANKING place="2" resultid="44" />
                    <RANKING place="1" resultid="1583" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2" agemax="11" agemin="10" name="Jahrgang 2012/2013">
                  <RANKINGS>
                    <RANKING place="2" resultid="582" />
                    <RANKING place="3" resultid="1573" />
                    <RANKING place="6" resultid="2167" />
                    <RANKING place="5" resultid="2177" />
                    <RANKING place="1" resultid="3978" />
                    <RANKING place="4" resultid="3981" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3" agemax="14" agemin="12" name="Jahrgang 2009 bis 2011">
                  <RANKINGS>
                    <RANKING place="6" resultid="28" />
                    <RANKING place="4" resultid="32" />
                    <RANKING place="15" resultid="575" />
                    <RANKING place="13" resultid="578" />
                    <RANKING place="8" resultid="602" />
                    <RANKING place="1" resultid="1536" />
                    <RANKING place="14" resultid="1551" />
                    <RANKING place="11" resultid="1555" />
                    <RANKING place="3" resultid="2149" />
                    <RANKING place="7" resultid="2160" />
                    <RANKING place="5" resultid="2179" />
                    <RANKING place="9" resultid="3987" />
                    <RANKING place="12" resultid="4010" />
                    <RANKING place="10" resultid="4016" />
                    <RANKING place="2" resultid="4183" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="17" agemin="15" name="Jahrgang 2006 bis 2008">
                  <RANKINGS>
                    <RANKING place="6" resultid="586" />
                    <RANKING place="10" resultid="598" />
                    <RANKING place="1" resultid="1559" />
                    <RANKING place="2" resultid="1577" />
                    <RANKING place="4" resultid="2169" />
                    <RANKING place="3" resultid="2173" />
                    <RANKING place="9" resultid="3993" />
                    <RANKING place="7" resultid="4000" />
                    <RANKING place="8" resultid="4004" />
                    <RANKING place="5" resultid="4019" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="50" number="112" gender="M" round="TIM">
              <SWIMSTYLE stroke="SURFACE" name="50 Flossenschwimmen Männer" relaycount="1" distance="50" />
              <HEATS>
                <HEAT heatid="50001" number="1" />
                <HEAT heatid="50002" number="2" />
                <HEAT heatid="50003" number="3" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="9" agemin="8" name="Jahrgang 2014/2015">
                  <RANKINGS>
                    <RANKING place="3" resultid="40" />
                    <RANKING place="2" resultid="48" />
                    <RANKING place="1" resultid="590" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2" agemax="11" agemin="10" name="Jahrgang 2012/2013">
                  <RANKINGS>
                    <RANKING place="4" resultid="568" />
                    <RANKING place="5" resultid="572" />
                    <RANKING place="3" resultid="594" />
                    <RANKING place="6" resultid="609" />
                    <RANKING place="1" resultid="1547" />
                    <RANKING place="2" resultid="2154" />
                    <RANKING place="7" resultid="2187" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3" agemax="14" agemin="12" name="Jahrgang 2009 bis 2011">
                  <RANKINGS>
                    <RANKING place="1" resultid="2144" />
                    <RANKING place="2" resultid="2157" />
                    <RANKING place="5" resultid="2163" />
                    <RANKING place="3" resultid="3975" />
                    <RANKING place="4" resultid="4007" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="17" agemin="15" name="Jahrgang 2006 bis 2008">
                  <RANKINGS>
                    <RANKING place="2" resultid="605" />
                    <RANKING place="3" resultid="1569" />
                    <RANKING place="1" resultid="2183" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
          </EVENTS>
        </SESSION>
        <SESSION number="3" date="2023-07-02" daytime="09:00" officialmeeting="08:30" warmupfrom="08:00">
          <EVENTS>
            <EVENT eventid="17" number="17" gender="F" round="TIM">
              <SWIMSTYLE stroke="BACK" name="50 Rückenbeinbewegung Frauen" technique="KICK" relaycount="1" distance="50" />
              <HEATS>
                <HEAT heatid="17001" number="1" />
                <HEAT heatid="17002" number="2" />
                <HEAT heatid="17003" number="3" />
                <HEAT heatid="17004" number="4" />
                <HEAT heatid="17005" number="5" />
                <HEAT heatid="17006" number="6" />
                <HEAT heatid="17007" number="7" />
                <HEAT heatid="17008" number="8" />
                <HEAT heatid="17009" number="9" />
                <HEAT heatid="17010" number="10" />
                <HEAT heatid="17011" number="11" />
                <HEAT heatid="17012" number="12" />
                <HEAT heatid="17013" number="13" />
                <HEAT heatid="17014" number="14" />
                <HEAT heatid="17015" number="15" />
                <HEAT heatid="17016" number="16" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="10" agemax="8" agemin="8" name="Jahrgang 2015">
                  <RANKINGS>
                    <RANKING place="8" resultid="197" />
                    <RANKING place="25" resultid="868" />
                    <RANKING place="10" resultid="879" />
                    <RANKING place="24" resultid="1928" />
                    <RANKING place="17" resultid="1976" />
                    <RANKING place="22" resultid="1981" />
                    <RANKING place="6" resultid="2077" />
                    <RANKING place="27" resultid="2081" />
                    <RANKING place="30" resultid="4088" />
                    <RANKING place="5" resultid="4201" />
                    <RANKING place="15" resultid="4218" />
                    <RANKING place="1" resultid="4222" />
                    <RANKING place="12" resultid="4226" />
                    <RANKING place="3" resultid="4336" />
                    <RANKING place="16" resultid="4350" />
                    <RANKING place="7" resultid="4384" />
                    <RANKING place="18" resultid="4413" />
                    <RANKING place="13" resultid="4470" />
                    <RANKING place="20" resultid="4667" />
                    <RANKING place="14" resultid="5005" />
                    <RANKING place="32" resultid="5040" />
                    <RANKING place="28" resultid="5054" />
                    <RANKING place="33" resultid="5089" />
                    <RANKING place="31" resultid="5122" />
                    <RANKING place="4" resultid="5126" />
                    <RANKING place="21" resultid="5200" />
                    <RANKING place="34" resultid="5855" />
                    <RANKING place="2" resultid="5965" />
                    <RANKING place="9" resultid="6006" />
                    <RANKING place="29" resultid="6074" />
                    <RANKING place="11" resultid="6128" />
                    <RANKING place="26" resultid="6132" />
                    <RANKING place="23" resultid="6172" />
                    <RANKING place="19" resultid="6228" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9" agemax="9" agemin="9" name="Jahrgang 2014">
                  <RANKINGS>
                    <RANKING place="31" resultid="227" />
                    <RANKING place="36" resultid="839" />
                    <RANKING place="11" resultid="911" />
                    <RANKING place="2" resultid="966" />
                    <RANKING place="6" resultid="1638" />
                    <RANKING place="1" resultid="1643" />
                    <RANKING place="23" resultid="1663" />
                    <RANKING place="24" resultid="1909" />
                    <RANKING place="35" resultid="1943" />
                    <RANKING place="16" resultid="2017" />
                    <RANKING place="32" resultid="2072" />
                    <RANKING place="30" resultid="4137" />
                    <RANKING place="12" resultid="4273" />
                    <RANKING place="17" resultid="4304" />
                    <RANKING place="9" resultid="4326" />
                    <RANKING place="13" resultid="4331" />
                    <RANKING place="14" resultid="4459" />
                    <RANKING place="40" resultid="4643" />
                    <RANKING place="19" resultid="5100" />
                    <RANKING place="4" resultid="5212" />
                    <RANKING place="29" resultid="5396" />
                    <RANKING place="37" resultid="5446" />
                    <RANKING place="15" resultid="5481" />
                    <RANKING place="39" resultid="5506" />
                    <RANKING place="20" resultid="5531" />
                    <RANKING place="18" resultid="5551" />
                    <RANKING place="8" resultid="5594" />
                    <RANKING place="34" resultid="5630" />
                    <RANKING place="27" resultid="5753" />
                    <RANKING place="26" resultid="5862" />
                    <RANKING place="7" resultid="5905" />
                    <RANKING place="21" resultid="6054" />
                    <RANKING place="10" resultid="6058" />
                    <RANKING place="33" resultid="6084" />
                    <RANKING place="38" resultid="6093" />
                    <RANKING place="25" resultid="6143" />
                    <RANKING place="3" resultid="6149" />
                    <RANKING place="5" resultid="6192" />
                    <RANKING place="28" resultid="6212" />
                    <RANKING place="22" resultid="6288" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1" agemax="10" agemin="10" name="Jahrgang 2013">
                  <RANKINGS>
                    <RANKING place="3" resultid="473" />
                    <RANKING place="12" resultid="842" />
                    <RANKING place="5" resultid="888" />
                    <RANKING place="17" resultid="950" />
                    <RANKING place="2" resultid="1919" />
                    <RANKING place="14" resultid="3494" />
                    <RANKING place="19" resultid="4299" />
                    <RANKING place="9" resultid="4357" />
                    <RANKING place="6" resultid="4428" />
                    <RANKING place="13" resultid="4473" />
                    <RANKING place="16" resultid="4635" />
                    <RANKING place="1" resultid="5442" />
                    <RANKING place="20" resultid="5464" />
                    <RANKING place="11" resultid="5725" />
                    <RANKING place="18" resultid="5770" />
                    <RANKING place="15" resultid="5780" />
                    <RANKING place="8" resultid="5925" />
                    <RANKING place="10" resultid="6043" />
                    <RANKING place="7" resultid="6050" />
                    <RANKING place="4" resultid="6107" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2" agemax="11" agemin="11" name="Jahrgang 2012">
                  <RANKINGS>
                    <RANKING place="3" resultid="957" />
                    <RANKING place="5" resultid="1597" />
                    <RANKING place="11" resultid="1614" />
                    <RANKING place="13" resultid="1651" />
                    <RANKING place="4" resultid="4322" />
                    <RANKING place="8" resultid="4813" />
                    <RANKING place="10" resultid="5108" />
                    <RANKING place="6" resultid="5180" />
                    <RANKING place="1" resultid="5343" />
                    <RANKING place="14" resultid="5612" />
                    <RANKING place="16" resultid="5817" />
                    <RANKING place="17" resultid="5858" />
                    <RANKING place="12" resultid="5974" />
                    <RANKING place="2" resultid="6037" />
                    <RANKING place="15" resultid="6302" />
                    <RANKING place="7" resultid="6333" />
                    <RANKING place="9" resultid="6339" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="18" number="18" gender="M" round="TIM">
              <SWIMSTYLE stroke="BACK" name="50 Rückenbeinbewegung Männer" technique="KICK" relaycount="1" distance="50" />
              <HEATS>
                <HEAT heatid="18001" number="1" />
                <HEAT heatid="18002" number="2" />
                <HEAT heatid="18003" number="3" />
                <HEAT heatid="18004" number="4" />
                <HEAT heatid="18005" number="5" />
                <HEAT heatid="18006" number="6" />
                <HEAT heatid="18007" number="7" />
                <HEAT heatid="18008" number="8" />
                <HEAT heatid="18009" number="9" />
                <HEAT heatid="18010" number="10" />
                <HEAT heatid="18011" number="11" />
                <HEAT heatid="18012" number="12" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="10" agemax="8" agemin="8" name="Jahrgang 2015">
                  <RANKINGS>
                    <RANKING place="22" resultid="193" />
                    <RANKING place="12" resultid="204" />
                    <RANKING place="16" resultid="215" />
                    <RANKING place="24" resultid="834" />
                    <RANKING place="15" resultid="864" />
                    <RANKING place="26" resultid="940" />
                    <RANKING place="20" resultid="970" />
                    <RANKING place="25" resultid="1886" />
                    <RANKING place="19" resultid="1899" />
                    <RANKING place="13" resultid="4079" />
                    <RANKING place="11" resultid="4163" />
                    <RANKING place="3" resultid="4184" />
                    <RANKING place="2" resultid="4375" />
                    <RANKING place="5" resultid="4522" />
                    <RANKING place="7" resultid="4665" />
                    <RANKING place="4" resultid="4674" />
                    <RANKING place="8" resultid="4679" />
                    <RANKING place="14" resultid="5014" />
                    <RANKING place="1" resultid="5653" />
                    <RANKING place="17" resultid="5969" />
                    <RANKING place="21" resultid="5987" />
                    <RANKING place="9" resultid="5990" />
                    <RANKING place="10" resultid="6014" />
                    <RANKING place="18" resultid="6066" />
                    <RANKING place="6" resultid="6103" />
                    <RANKING place="23" resultid="6206" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9" agemax="9" agemin="9" name="Jahrgang 2014">
                  <RANKINGS>
                    <RANKING place="28" resultid="236" />
                    <RANKING place="1" resultid="884" />
                    <RANKING place="8" resultid="983" />
                    <RANKING place="19" resultid="1605" />
                    <RANKING place="17" resultid="1971" />
                    <RANKING place="7" resultid="2003" />
                    <RANKING place="32" resultid="2022" />
                    <RANKING place="25" resultid="2053" />
                    <RANKING place="22" resultid="4115" />
                    <RANKING place="16" resultid="4142" />
                    <RANKING place="27" resultid="4188" />
                    <RANKING place="5" resultid="4205" />
                    <RANKING place="33" resultid="4209" />
                    <RANKING place="4" resultid="4230" />
                    <RANKING place="15" resultid="4235" />
                    <RANKING place="11" resultid="4532" />
                    <RANKING place="24" resultid="4769" />
                    <RANKING place="26" resultid="5183" />
                    <RANKING place="30" resultid="5195" />
                    <RANKING place="9" resultid="5467" />
                    <RANKING place="3" resultid="5599" />
                    <RANKING place="14" resultid="5692" />
                    <RANKING place="2" resultid="5904" />
                    <RANKING place="20" resultid="5957" />
                    <RANKING place="12" resultid="5994" />
                    <RANKING place="13" resultid="6153" />
                    <RANKING place="6" resultid="6216" />
                    <RANKING place="18" resultid="6238" />
                    <RANKING place="10" resultid="6241" />
                    <RANKING place="31" resultid="6254" />
                    <RANKING place="21" resultid="6278" />
                    <RANKING place="29" resultid="6353" />
                    <RANKING place="23" resultid="6356" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1" agemax="10" agemin="10" name="Jahrgang 2013">
                  <RANKINGS>
                    <RANKING place="6" resultid="2131" />
                    <RANKING place="10" resultid="3738" />
                    <RANKING place="5" resultid="4421" />
                    <RANKING place="3" resultid="4497" />
                    <RANKING place="2" resultid="5538" />
                    <RANKING place="9" resultid="5542" />
                    <RANKING place="4" resultid="5837" />
                    <RANKING place="1" resultid="5889" />
                    <RANKING place="8" resultid="6266" />
                    <RANKING place="7" resultid="6312" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2" agemax="11" agemin="11" name="Jahrgang 2012">
                  <RANKINGS>
                    <RANKING place="1" resultid="125" />
                    <RANKING place="7" resultid="201" />
                    <RANKING place="11" resultid="813" />
                    <RANKING place="12" resultid="857" />
                    <RANKING place="10" resultid="991" />
                    <RANKING place="9" resultid="4269" />
                    <RANKING place="6" resultid="4348" />
                    <RANKING place="4" resultid="4451" />
                    <RANKING place="2" resultid="5527" />
                    <RANKING place="8" resultid="5568" />
                    <RANKING place="5" resultid="5804" />
                    <RANKING place="15" resultid="5810" />
                    <RANKING place="3" resultid="5851" />
                    <RANKING place="13" resultid="6269" />
                    <RANKING place="14" resultid="6299" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="19" number="19" gender="F" round="TIM">
              <SWIMSTYLE stroke="BREAST" relaycount="1" distance="50" />
              <HEATS>
                <HEAT heatid="19001" number="1" />
                <HEAT heatid="19002" number="2" />
                <HEAT heatid="19003" number="3" />
                <HEAT heatid="19004" number="4" />
                <HEAT heatid="19005" number="5" />
                <HEAT heatid="19006" number="6" />
                <HEAT heatid="19007" number="7" />
                <HEAT heatid="19008" number="8" />
                <HEAT heatid="19009" number="9" />
                <HEAT heatid="19010" number="10" />
                <HEAT heatid="19011" number="11" />
                <HEAT heatid="19012" number="12" />
                <HEAT heatid="19013" number="13" />
                <HEAT heatid="19014" number="14" />
                <HEAT heatid="19015" number="15" />
                <HEAT heatid="19016" number="16" />
                <HEAT heatid="19017" number="17" />
                <HEAT heatid="19018" number="18" />
                <HEAT heatid="19019" number="19" />
                <HEAT heatid="19020" number="20" />
                <HEAT heatid="19021" number="21" />
                <HEAT heatid="19022" number="22" />
                <HEAT heatid="19023" number="23" />
                <HEAT heatid="19024" number="24" />
                <HEAT heatid="19025" number="25" />
                <HEAT heatid="19026" number="26" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="10" agemax="8" agemin="8" name="Jahrgang 2015">
                  <RANKINGS>
                    <RANKING place="16" resultid="220" />
                    <RANKING place="26" resultid="902" />
                    <RANKING place="20" resultid="906" />
                    <RANKING place="21" resultid="1006" />
                    <RANKING place="13" resultid="1903" />
                    <RANKING place="33" resultid="1927" />
                    <RANKING place="31" resultid="1975" />
                    <RANKING place="25" resultid="1980" />
                    <RANKING place="29" resultid="2076" />
                    <RANKING place="4" resultid="3449" />
                    <RANKING place="7" resultid="3832" />
                    <RANKING place="38" resultid="4055" />
                    <RANKING place="30" resultid="4251" />
                    <RANKING place="3" resultid="4340" />
                    <RANKING place="11" resultid="4425" />
                    <RANKING place="9" resultid="4448" />
                    <RANKING place="27" resultid="4485" />
                    <RANKING place="6" resultid="4489" />
                    <RANKING place="14" resultid="4526" />
                    <RANKING place="5" resultid="4585" />
                    <RANKING place="28" resultid="4937" />
                    <RANKING place="39" resultid="5006" />
                    <RANKING place="40" resultid="5055" />
                    <RANKING place="24" resultid="5072" />
                    <RANKING place="15" resultid="5090" />
                    <RANKING place="17" resultid="5118" />
                    <RANKING place="35" resultid="5123" />
                    <RANKING place="10" resultid="5127" />
                    <RANKING place="8" resultid="5201" />
                    <RANKING place="22" resultid="5224" />
                    <RANKING place="23" resultid="5856" />
                    <RANKING place="1" resultid="5966" />
                    <RANKING place="18" resultid="5980" />
                    <RANKING place="12" resultid="6007" />
                    <RANKING place="34" resultid="6090" />
                    <RANKING place="19" resultid="6111" />
                    <RANKING place="32" resultid="6133" />
                    <RANKING place="36" resultid="6173" />
                    <RANKING place="37" resultid="6229" />
                    <RANKING place="2" resultid="6295" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9" agemax="9" agemin="9" name="Jahrgang 2014">
                  <RANKINGS>
                    <RANKING place="2" resultid="803" />
                    <RANKING place="17" resultid="923" />
                    <RANKING place="19" resultid="936" />
                    <RANKING place="12" resultid="1637" />
                    <RANKING place="29" resultid="1658" />
                    <RANKING place="14" resultid="1908" />
                    <RANKING place="45" resultid="1942" />
                    <RANKING place="41" resultid="2071" />
                    <RANKING place="25" resultid="2097" />
                    <RANKING place="6" resultid="3480" />
                    <RANKING place="42" resultid="3719" />
                    <RANKING place="32" resultid="4083" />
                    <RANKING place="46" resultid="4093" />
                    <RANKING place="24" resultid="4120" />
                    <RANKING place="44" resultid="4138" />
                    <RANKING place="43" resultid="4148" />
                    <RANKING place="1" resultid="4278" />
                    <RANKING place="9" resultid="4309" />
                    <RANKING place="21" resultid="4361" />
                    <RANKING place="36" resultid="4370" />
                    <RANKING place="7" resultid="4380" />
                    <RANKING place="3" resultid="4408" />
                    <RANKING place="16" resultid="4432" />
                    <RANKING place="38" resultid="5019" />
                    <RANKING place="40" resultid="5024" />
                    <RANKING place="22" resultid="5044" />
                    <RANKING place="37" resultid="5101" />
                    <RANKING place="11" resultid="5112" />
                    <RANKING place="27" resultid="5290" />
                    <RANKING place="5" resultid="5376" />
                    <RANKING place="13" resultid="5380" />
                    <RANKING place="28" resultid="5397" />
                    <RANKING place="10" resultid="5447" />
                    <RANKING place="23" resultid="5482" />
                    <RANKING place="33" resultid="5507" />
                    <RANKING place="31" resultid="5532" />
                    <RANKING place="34" resultid="5552" />
                    <RANKING place="8" resultid="5631" />
                    <RANKING place="4" resultid="5676" />
                    <RANKING place="20" resultid="5754" />
                    <RANKING place="25" resultid="5864" />
                    <RANKING place="39" resultid="5868" />
                    <RANKING place="15" resultid="6055" />
                    <RANKING place="48" resultid="6085" />
                    <RANKING place="47" resultid="6094" />
                    <RANKING place="18" resultid="6144" />
                    <RANKING place="35" resultid="6150" />
                    <RANKING place="30" resultid="6193" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1" agemax="10" agemin="10" name="Jahrgang 2013">
                  <RANKINGS>
                    <RANKING place="5" resultid="211" />
                    <RANKING place="14" resultid="245" />
                    <RANKING place="13" resultid="763" />
                    <RANKING place="4" resultid="766" />
                    <RANKING place="9" resultid="781" />
                    <RANKING place="8" resultid="799" />
                    <RANKING place="25" resultid="1966" />
                    <RANKING place="10" resultid="1998" />
                    <RANKING place="15" resultid="3826" />
                    <RANKING place="23" resultid="4128" />
                    <RANKING place="24" resultid="4160" />
                    <RANKING place="18" resultid="4353" />
                    <RANKING place="3" resultid="4444" />
                    <RANKING place="2" resultid="4455" />
                    <RANKING place="16" resultid="4617" />
                    <RANKING place="19" resultid="4636" />
                    <RANKING place="6" resultid="4749" />
                    <RANKING place="12" resultid="5096" />
                    <RANKING place="1" resultid="5221" />
                    <RANKING place="20" resultid="5465" />
                    <RANKING place="11" resultid="5477" />
                    <RANKING place="26" resultid="5726" />
                    <RANKING place="22" resultid="5781" />
                    <RANKING place="7" resultid="5831" />
                    <RANKING place="17" resultid="5926" />
                    <RANKING place="21" resultid="6324" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2" agemax="11" agemin="11" name="Jahrgang 2012">
                  <RANKINGS>
                    <RANKING place="8" resultid="181" />
                    <RANKING place="2" resultid="1893" />
                    <RANKING place="6" resultid="1951" />
                    <RANKING place="20" resultid="3812" />
                    <RANKING place="1" resultid="4438" />
                    <RANKING place="19" resultid="4477" />
                    <RANKING place="25" resultid="4561" />
                    <RANKING place="11" resultid="4814" />
                    <RANKING place="12" resultid="4859" />
                    <RANKING place="18" resultid="4874" />
                    <RANKING place="22" resultid="4920" />
                    <RANKING place="16" resultid="5036" />
                    <RANKING place="10" resultid="5232" />
                    <RANKING place="9" resultid="5493" />
                    <RANKING place="20" resultid="5619" />
                    <RANKING place="3" resultid="5638" />
                    <RANKING place="7" resultid="5645" />
                    <RANKING place="24" resultid="5672" />
                    <RANKING place="5" resultid="5713" />
                    <RANKING place="14" resultid="5721" />
                    <RANKING place="17" resultid="5859" />
                    <RANKING place="13" resultid="6025" />
                    <RANKING place="15" resultid="6179" />
                    <RANKING place="23" resultid="6303" />
                    <RANKING place="4" resultid="6347" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="13" agemin="12" name="Jahrgang 2010/2011">
                  <RANKINGS>
                    <RANKING place="1" resultid="133" />
                    <RANKING place="3" resultid="149" />
                    <RANKING place="12" resultid="157" />
                    <RANKING place="4" resultid="173" />
                    <RANKING place="31" resultid="224" />
                    <RANKING place="18" resultid="1987" />
                    <RANKING place="21" resultid="2061" />
                    <RANKING place="32" resultid="2101" />
                    <RANKING place="28" resultid="2105" />
                    <RANKING place="2" resultid="2139" />
                    <RANKING place="16" resultid="3760" />
                    <RANKING place="34" resultid="3780" />
                    <RANKING place="30" resultid="4301" />
                    <RANKING place="10" resultid="4442" />
                    <RANKING place="9" resultid="4548" />
                    <RANKING place="33" resultid="4559" />
                    <RANKING place="26" resultid="4697" />
                    <RANKING place="17" resultid="4846" />
                    <RANKING place="15" resultid="4867" />
                    <RANKING place="7" resultid="4881" />
                    <RANKING place="25" resultid="5002" />
                    <RANKING place="23" resultid="5029" />
                    <RANKING place="22" resultid="5086" />
                    <RANKING place="13" resultid="5148" />
                    <RANKING place="5" resultid="5209" />
                    <RANKING place="27" resultid="5370" />
                    <RANKING place="6" resultid="5404" />
                    <RANKING place="29" resultid="5504" />
                    <RANKING place="19" resultid="5549" />
                    <RANKING place="24" resultid="5762" />
                    <RANKING place="14" resultid="5777" />
                    <RANKING place="20" resultid="5790" />
                    <RANKING place="11" resultid="6285" />
                    <RANKING place="8" resultid="6360" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6" agemax="15" agemin="14" name="Jahrgang 2008/2009">
                  <RANKINGS>
                    <RANKING place="14" resultid="3461" />
                    <RANKING place="2" resultid="3821" />
                    <RANKING place="11" resultid="4290" />
                    <RANKING place="1" resultid="4581" />
                    <RANKING place="13" resultid="4744" />
                    <RANKING place="5" resultid="4887" />
                    <RANKING place="6" resultid="4943" />
                    <RANKING place="8" resultid="4978" />
                    <RANKING place="15" resultid="5294" />
                    <RANKING place="3" resultid="5498" />
                    <RANKING place="4" resultid="5651" />
                    <RANKING place="9" resultid="5921" />
                    <RANKING place="7" resultid="5963" />
                    <RANKING place="12" resultid="6158" />
                    <RANKING place="10" resultid="6190" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8" agemax="17" agemin="16" name="Jahrgang 2006/2007">
                  <RANKINGS>
                    <RANKING place="2" resultid="4651" />
                    <RANKING place="1" resultid="4840" />
                    <RANKING place="3" resultid="4960" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="20" number="20" gender="M" round="TIM">
              <SWIMSTYLE stroke="BREAST" relaycount="1" distance="50" />
              <HEATS>
                <HEAT heatid="20001" number="1" />
                <HEAT heatid="20002" number="2" />
                <HEAT heatid="20003" number="3" />
                <HEAT heatid="20004" number="4" />
                <HEAT heatid="20005" number="5" />
                <HEAT heatid="20006" number="6" />
                <HEAT heatid="20007" number="7" />
                <HEAT heatid="20008" number="8" />
                <HEAT heatid="20009" number="9" />
                <HEAT heatid="20010" number="10" />
                <HEAT heatid="20011" number="11" />
                <HEAT heatid="20012" number="12" />
                <HEAT heatid="20013" number="13" />
                <HEAT heatid="20014" number="14" />
                <HEAT heatid="20015" number="15" />
                <HEAT heatid="20016" number="16" />
                <HEAT heatid="20017" number="17" />
                <HEAT heatid="20018" number="18" />
                <HEAT heatid="20019" number="19" />
                <HEAT heatid="20020" number="20" />
                <HEAT heatid="20021" number="21" />
                <HEAT heatid="20022" number="22" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="10" agemax="8" agemin="8" name="Jahrgang 2015">
                  <RANKINGS>
                    <RANKING place="17" resultid="863" />
                    <RANKING place="20" resultid="931" />
                    <RANKING place="6" resultid="1898" />
                    <RANKING place="7" resultid="2030" />
                    <RANKING place="23" resultid="2067" />
                    <RANKING place="1" resultid="3844" />
                    <RANKING place="19" resultid="4080" />
                    <RANKING place="9" resultid="4376" />
                    <RANKING place="2" resultid="4396" />
                    <RANKING place="8" resultid="4493" />
                    <RANKING place="4" resultid="4518" />
                    <RANKING place="3" resultid="4675" />
                    <RANKING place="24" resultid="4712" />
                    <RANKING place="22" resultid="4788" />
                    <RANKING place="11" resultid="5015" />
                    <RANKING place="5" resultid="5654" />
                    <RANKING place="25" resultid="5970" />
                    <RANKING place="21" resultid="5984" />
                    <RANKING place="18" resultid="5991" />
                    <RANKING place="16" resultid="6067" />
                    <RANKING place="15" resultid="6071" />
                    <RANKING place="10" resultid="6122" />
                    <RANKING place="12" resultid="6163" />
                    <RANKING place="13" resultid="6203" />
                    <RANKING place="14" resultid="6225" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9" agemax="9" agemin="9" name="Jahrgang 2014">
                  <RANKINGS>
                    <RANKING place="15" resultid="477" />
                    <RANKING place="17" resultid="927" />
                    <RANKING place="25" resultid="987" />
                    <RANKING place="28" resultid="1010" />
                    <RANKING place="7" resultid="1020" />
                    <RANKING place="2" resultid="1621" />
                    <RANKING place="19" resultid="1970" />
                    <RANKING place="29" resultid="2021" />
                    <RANKING place="30" resultid="2052" />
                    <RANKING place="3" resultid="2058" />
                    <RANKING place="6" resultid="4024" />
                    <RANKING place="13" resultid="4032" />
                    <RANKING place="8" resultid="4045" />
                    <RANKING place="26" resultid="4116" />
                    <RANKING place="5" resultid="4189" />
                    <RANKING place="10" resultid="4192" />
                    <RANKING place="12" resultid="4196" />
                    <RANKING place="1" resultid="4210" />
                    <RANKING place="23" resultid="4236" />
                    <RANKING place="22" resultid="4533" />
                    <RANKING place="16" resultid="4654" />
                    <RANKING place="27" resultid="5184" />
                    <RANKING place="31" resultid="5196" />
                    <RANKING place="9" resultid="5407" />
                    <RANKING place="11" resultid="5693" />
                    <RANKING place="4" resultid="5728" />
                    <RANKING place="20" resultid="5995" />
                    <RANKING place="18" resultid="6217" />
                    <RANKING place="21" resultid="6239" />
                    <RANKING place="14" resultid="6255" />
                    <RANKING place="32" resultid="6342" />
                    <RANKING place="24" resultid="6354" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1" agemax="10" agemin="10" name="Jahrgang 2013">
                  <RANKINGS>
                    <RANKING place="7" resultid="760" />
                    <RANKING place="5" resultid="850" />
                    <RANKING place="14" resultid="1624" />
                    <RANKING place="6" resultid="1630" />
                    <RANKING place="21" resultid="2037" />
                    <RANKING place="17" resultid="3497" />
                    <RANKING place="16" resultid="3840" />
                    <RANKING place="3" resultid="4041" />
                    <RANKING place="11" resultid="4052" />
                    <RANKING place="9" resultid="4100" />
                    <RANKING place="19" resultid="4249" />
                    <RANKING place="15" resultid="4344" />
                    <RANKING place="2" resultid="4366" />
                    <RANKING place="8" resultid="4761" />
                    <RANKING place="18" resultid="5064" />
                    <RANKING place="22" resultid="5543" />
                    <RANKING place="1" resultid="5588" />
                    <RANKING place="12" resultid="5945" />
                    <RANKING place="4" resultid="5953" />
                    <RANKING place="10" resultid="6199" />
                    <RANKING place="13" resultid="6262" />
                    <RANKING place="20" resultid="6313" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2" agemax="11" agemin="11" name="Jahrgang 2012">
                  <RANKINGS>
                    <RANKING place="20" resultid="202" />
                    <RANKING place="13" resultid="784" />
                    <RANKING place="4" resultid="820" />
                    <RANKING place="5" resultid="2007" />
                    <RANKING place="1" resultid="3457" />
                    <RANKING place="17" resultid="3749" />
                    <RANKING place="15" resultid="3789" />
                    <RANKING place="8" resultid="4067" />
                    <RANKING place="19" resultid="4170" />
                    <RANKING place="3" resultid="4400" />
                    <RANKING place="12" resultid="4719" />
                    <RANKING place="6" resultid="4726" />
                    <RANKING place="9" resultid="4827" />
                    <RANKING place="7" resultid="5309" />
                    <RANKING place="2" resultid="5519" />
                    <RANKING place="14" resultid="5805" />
                    <RANKING place="18" resultid="5811" />
                    <RANKING place="10" resultid="6010" />
                    <RANKING place="11" resultid="6252" />
                    <RANKING place="16" resultid="6270" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="13" agemin="12" name="Jahrgang 2010/2011">
                  <RANKINGS>
                    <RANKING place="8" resultid="117" />
                    <RANKING place="6" resultid="141" />
                    <RANKING place="2" resultid="770" />
                    <RANKING place="9" resultid="792" />
                    <RANKING place="7" resultid="810" />
                    <RANKING place="5" resultid="871" />
                    <RANKING place="30" resultid="1890" />
                    <RANKING place="24" resultid="1931" />
                    <RANKING place="18" resultid="2048" />
                    <RANKING place="29" resultid="2090" />
                    <RANKING place="4" resultid="3442" />
                    <RANKING place="20" resultid="3734" />
                    <RANKING place="32" resultid="3848" />
                    <RANKING place="12" resultid="4287" />
                    <RANKING place="3" resultid="4468" />
                    <RANKING place="10" resultid="4554" />
                    <RANKING place="19" resultid="4571" />
                    <RANKING place="11" resultid="4593" />
                    <RANKING place="1" resultid="4629" />
                    <RANKING place="31" resultid="4641" />
                    <RANKING place="22" resultid="4893" />
                    <RANKING place="26" resultid="4901" />
                    <RANKING place="23" resultid="4988" />
                    <RANKING place="13" resultid="5243" />
                    <RANKING place="16" resultid="5426" />
                    <RANKING place="25" resultid="5512" />
                    <RANKING place="21" resultid="5661" />
                    <RANKING place="14" resultid="5749" />
                    <RANKING place="15" resultid="5883" />
                    <RANKING place="17" resultid="6166" />
                    <RANKING place="26" resultid="6309" />
                    <RANKING place="28" resultid="6330" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6" agemax="15" agemin="14" name="Jahrgang 2008/2009">
                  <RANKINGS>
                    <RANKING place="16" resultid="3491" />
                    <RANKING place="9" resultid="3714" />
                    <RANKING place="2" resultid="3775" />
                    <RANKING place="6" resultid="3817" />
                    <RANKING place="12" resultid="4263" />
                    <RANKING place="1" resultid="4317" />
                    <RANKING place="18" resultid="4538" />
                    <RANKING place="13" resultid="4600" />
                    <RANKING place="11" resultid="4662" />
                    <RANKING place="19" resultid="4807" />
                    <RANKING place="17" resultid="4821" />
                    <RANKING place="7" resultid="4853" />
                    <RANKING place="15" resultid="4907" />
                    <RANKING place="3" resultid="4953" />
                    <RANKING place="10" resultid="5068" />
                    <RANKING place="4" resultid="5362" />
                    <RANKING place="5" resultid="5768" />
                    <RANKING place="8" resultid="6082" />
                    <RANKING place="14" resultid="6097" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8" agemax="17" agemin="16" name="Jahrgang 2006/2007">
                  <RANKINGS>
                    <RANKING place="1" resultid="3465" />
                    <RANKING place="5" resultid="3484" />
                    <RANKING place="8" resultid="3797" />
                    <RANKING place="7" resultid="4297" />
                    <RANKING place="9" resultid="4834" />
                    <RANKING place="2" resultid="5135" />
                    <RANKING place="4" resultid="5372" />
                    <RANKING place="3" resultid="5582" />
                    <RANKING place="6" resultid="6306" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="21" number="21" gender="F" round="TIM">
              <SWIMSTYLE stroke="FREE" name="50 Kraulbeinbewegung Frauen" technique="KICK" relaycount="1" distance="50" />
              <HEATS>
                <HEAT heatid="21001" number="1" />
                <HEAT heatid="21002" number="2" />
                <HEAT heatid="21003" number="3" />
                <HEAT heatid="21004" number="4" />
                <HEAT heatid="21005" number="5" />
                <HEAT heatid="21006" number="6" />
                <HEAT heatid="21007" number="7" />
                <HEAT heatid="21008" number="8" />
                <HEAT heatid="21009" number="9" />
                <HEAT heatid="21010" number="10" />
                <HEAT heatid="21011" number="11" />
                <HEAT heatid="21012" number="12" />
                <HEAT heatid="21013" number="13" />
                <HEAT heatid="21014" number="14" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="10" agemax="8" agemin="8" name="Jahrgang 2015">
                  <RANKINGS>
                    <RANKING place="11" resultid="198" />
                    <RANKING place="28" resultid="221" />
                    <RANKING place="29" resultid="867" />
                    <RANKING place="4" resultid="878" />
                    <RANKING place="22" resultid="1902" />
                    <RANKING place="8" resultid="1974" />
                    <RANKING place="32" resultid="2080" />
                    <RANKING place="27" resultid="4056" />
                    <RANKING place="21" resultid="4089" />
                    <RANKING place="19" resultid="4154" />
                    <RANKING place="1" resultid="4202" />
                    <RANKING place="15" resultid="4219" />
                    <RANKING place="13" resultid="4223" />
                    <RANKING place="6" resultid="4227" />
                    <RANKING place="19" resultid="4252" />
                    <RANKING place="3" resultid="4337" />
                    <RANKING place="2" resultid="4341" />
                    <RANKING place="14" resultid="4351" />
                    <RANKING place="9" resultid="4385" />
                    <RANKING place="25" resultid="4414" />
                    <RANKING place="12" resultid="4471" />
                    <RANKING place="24" resultid="4486" />
                    <RANKING place="18" resultid="4586" />
                    <RANKING place="26" resultid="4668" />
                    <RANKING place="31" resultid="5041" />
                    <RANKING place="33" resultid="5073" />
                    <RANKING place="23" resultid="5091" />
                    <RANKING place="16" resultid="5225" />
                    <RANKING place="10" resultid="5981" />
                    <RANKING place="17" resultid="6008" />
                    <RANKING place="30" resultid="6075" />
                    <RANKING place="7" resultid="6129" />
                    <RANKING place="5" resultid="6296" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9" agemax="9" agemin="9" name="Jahrgang 2014">
                  <RANKINGS>
                    <RANKING place="32" resultid="228" />
                    <RANKING place="33" resultid="838" />
                    <RANKING place="19" resultid="922" />
                    <RANKING place="1" resultid="1642" />
                    <RANKING place="28" resultid="1662" />
                    <RANKING place="30" resultid="2016" />
                    <RANKING place="31" resultid="2070" />
                    <RANKING place="16" resultid="2096" />
                    <RANKING place="21" resultid="3452" />
                    <RANKING place="2" resultid="4121" />
                    <RANKING place="11" resultid="4139" />
                    <RANKING place="3" resultid="4274" />
                    <RANKING place="23" resultid="4305" />
                    <RANKING place="8" resultid="4327" />
                    <RANKING place="20" resultid="4332" />
                    <RANKING place="26" resultid="4362" />
                    <RANKING place="9" resultid="4371" />
                    <RANKING place="24" resultid="4409" />
                    <RANKING place="5" resultid="4765" />
                    <RANKING place="22" resultid="5025" />
                    <RANKING place="25" resultid="5077" />
                    <RANKING place="15" resultid="5213" />
                    <RANKING place="29" resultid="5291" />
                    <RANKING place="7" resultid="5381" />
                    <RANKING place="10" resultid="5559" />
                    <RANKING place="12" resultid="5595" />
                    <RANKING place="6" resultid="5677" />
                    <RANKING place="13" resultid="5755" />
                    <RANKING place="4" resultid="5865" />
                    <RANKING place="17" resultid="5906" />
                    <RANKING place="18" resultid="6059" />
                    <RANKING place="14" resultid="6213" />
                    <RANKING place="27" resultid="6289" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1" agemax="10" agemin="10" name="Jahrgang 2013">
                  <RANKINGS>
                    <RANKING place="11" resultid="841" />
                    <RANKING place="6" resultid="887" />
                    <RANKING place="14" resultid="949" />
                    <RANKING place="21" resultid="1965" />
                    <RANKING place="15" resultid="3493" />
                    <RANKING place="12" resultid="3729" />
                    <RANKING place="18" resultid="4129" />
                    <RANKING place="20" resultid="4161" />
                    <RANKING place="16" resultid="4300" />
                    <RANKING place="2" resultid="4429" />
                    <RANKING place="7" resultid="4510" />
                    <RANKING place="5" resultid="4514" />
                    <RANKING place="10" resultid="4618" />
                    <RANKING place="8" resultid="4692" />
                    <RANKING place="1" resultid="5142" />
                    <RANKING place="3" resultid="5222" />
                    <RANKING place="4" resultid="5576" />
                    <RANKING place="19" resultid="5727" />
                    <RANKING place="17" resultid="5771" />
                    <RANKING place="13" resultid="6044" />
                    <RANKING place="9" resultid="6051" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2" agemax="11" agemin="11" name="Jahrgang 2012">
                  <RANKINGS>
                    <RANKING place="4" resultid="1608" />
                    <RANKING place="8" resultid="1646" />
                    <RANKING place="2" resultid="4323" />
                    <RANKING place="6" resultid="4913" />
                    <RANKING place="1" resultid="5181" />
                    <RANKING place="7" resultid="5620" />
                    <RANKING place="11" resultid="5818" />
                    <RANKING place="3" resultid="5933" />
                    <RANKING place="9" resultid="6026" />
                    <RANKING place="5" resultid="6334" />
                    <RANKING place="10" resultid="6340" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="22" number="22" gender="M" round="TIM">
              <SWIMSTYLE stroke="FREE" name="50 Kraulbeinbewegung Männer" technique="KICK" relaycount="1" distance="50" />
              <HEATS>
                <HEAT heatid="22001" number="1" />
                <HEAT heatid="22002" number="2" />
                <HEAT heatid="22003" number="3" />
                <HEAT heatid="22004" number="4" />
                <HEAT heatid="22005" number="5" />
                <HEAT heatid="22006" number="6" />
                <HEAT heatid="22007" number="7" />
                <HEAT heatid="22008" number="8" />
                <HEAT heatid="22009" number="9" />
                <HEAT heatid="22010" number="10" />
                <HEAT heatid="22011" number="11" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="10" agemax="8" agemin="8" name="Jahrgang 2015">
                  <RANKINGS>
                    <RANKING place="16" resultid="194" />
                    <RANKING place="7" resultid="205" />
                    <RANKING place="17" resultid="216" />
                    <RANKING place="6" resultid="939" />
                    <RANKING place="11" resultid="969" />
                    <RANKING place="22" resultid="1885" />
                    <RANKING place="14" resultid="3843" />
                    <RANKING place="3" resultid="4164" />
                    <RANKING place="2" resultid="4185" />
                    <RANKING place="1" resultid="4377" />
                    <RANKING place="12" resultid="4397" />
                    <RANKING place="5" resultid="4523" />
                    <RANKING place="9" resultid="4666" />
                    <RANKING place="4" resultid="4676" />
                    <RANKING place="10" resultid="4680" />
                    <RANKING place="20" resultid="4713" />
                    <RANKING place="21" resultid="5016" />
                    <RANKING place="18" resultid="5988" />
                    <RANKING place="15" resultid="5992" />
                    <RANKING place="8" resultid="6015" />
                    <RANKING place="23" resultid="6204" />
                    <RANKING place="13" resultid="6207" />
                    <RANKING place="19" resultid="6226" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9" agemax="9" agemin="9" name="Jahrgang 2014">
                  <RANKINGS>
                    <RANKING place="25" resultid="237" />
                    <RANKING place="14" resultid="478" />
                    <RANKING place="1" resultid="883" />
                    <RANKING place="10" resultid="1604" />
                    <RANKING place="6" resultid="2002" />
                    <RANKING place="28" resultid="2020" />
                    <RANKING place="23" resultid="2051" />
                    <RANKING place="5" resultid="2057" />
                    <RANKING place="27" resultid="4033" />
                    <RANKING place="15" resultid="4046" />
                    <RANKING place="22" resultid="4117" />
                    <RANKING place="4" resultid="4143" />
                    <RANKING place="17" resultid="4190" />
                    <RANKING place="11" resultid="4197" />
                    <RANKING place="7" resultid="4206" />
                    <RANKING place="12" resultid="4237" />
                    <RANKING place="18" resultid="4770" />
                    <RANKING place="16" resultid="5049" />
                    <RANKING place="3" resultid="5600" />
                    <RANKING place="13" resultid="5694" />
                    <RANKING place="2" resultid="5729" />
                    <RANKING place="24" resultid="5958" />
                    <RANKING place="20" resultid="5996" />
                    <RANKING place="19" resultid="6154" />
                    <RANKING place="9" resultid="6240" />
                    <RANKING place="8" resultid="6242" />
                    <RANKING place="21" resultid="6279" />
                    <RANKING place="26" resultid="6357" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1" agemax="10" agemin="10" name="Jahrgang 2013">
                  <RANKINGS>
                    <RANKING place="4" resultid="1623" />
                    <RANKING place="11" resultid="2036" />
                    <RANKING place="1" resultid="3436" />
                    <RANKING place="10" resultid="3737" />
                    <RANKING place="8" resultid="3839" />
                    <RANKING place="7" resultid="4392" />
                    <RANKING place="9" resultid="4778" />
                    <RANKING place="2" resultid="4984" />
                    <RANKING place="5" resultid="5173" />
                    <RANKING place="3" resultid="5626" />
                    <RANKING place="6" resultid="5890" />
                    <RANKING place="12" resultid="6267" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2" agemax="11" agemin="11" name="Jahrgang 2012">
                  <RANKINGS>
                    <RANKING place="1" resultid="189" />
                    <RANKING place="8" resultid="999" />
                    <RANKING place="4" resultid="2135" />
                    <RANKING place="13" resultid="3748" />
                    <RANKING place="11" resultid="4171" />
                    <RANKING place="2" resultid="4242" />
                    <RANKING place="6" resultid="4270" />
                    <RANKING place="3" resultid="4417" />
                    <RANKING place="10" resultid="4481" />
                    <RANKING place="5" resultid="4798" />
                    <RANKING place="9" resultid="5569" />
                    <RANKING place="7" resultid="5852" />
                    <RANKING place="12" resultid="6271" />
                    <RANKING place="14" resultid="6300" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="23" number="23" gender="F" round="TIM">
              <SWIMSTYLE stroke="FREE" relaycount="1" distance="200" />
              <HEATS>
                <HEAT heatid="23001" number="1" />
                <HEAT heatid="23002" number="2" />
                <HEAT heatid="23003" number="3" />
                <HEAT heatid="23004" number="4" />
                <HEAT heatid="23005" number="5" />
                <HEAT heatid="23006" number="6" />
                <HEAT heatid="23007" number="7" />
                <HEAT heatid="23008" number="8" />
                <HEAT heatid="23009" number="9" />
                <HEAT heatid="23010" number="10" />
                <HEAT heatid="23011" number="11" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="10" agemin="10" name="Jahrgang 2013">
                  <RANKINGS>
                    <RANKING place="4" resultid="212" />
                    <RANKING place="3" resultid="246" />
                    <RANKING place="6" resultid="840" />
                    <RANKING place="10" resultid="4354" />
                    <RANKING place="1" resultid="4511" />
                    <RANKING place="2" resultid="4515" />
                    <RANKING place="8" resultid="4693" />
                    <RANKING place="7" resultid="5192" />
                    <RANKING place="9" resultid="5478" />
                    <RANKING place="5" resultid="5577" />
                    <RANKING place="11" resultid="5927" />
                    <RANKING place="12" resultid="6045" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2" agemax="11" agemin="11" name="Jahrgang 2012">
                  <RANKINGS>
                    <RANKING place="5" resultid="18" />
                    <RANKING place="12" resultid="1613" />
                    <RANKING place="15" resultid="1650" />
                    <RANKING place="14" resultid="1892" />
                    <RANKING place="17" resultid="1950" />
                    <RANKING place="2" resultid="1955" />
                    <RANKING place="7" resultid="1992" />
                    <RANKING place="1" resultid="4439" />
                    <RANKING place="10" resultid="4478" />
                    <RANKING place="9" resultid="4503" />
                    <RANKING place="4" resultid="4507" />
                    <RANKING place="3" resultid="4740" />
                    <RANKING place="16" resultid="5613" />
                    <RANKING place="8" resultid="5844" />
                    <RANKING place="13" resultid="5934" />
                    <RANKING place="11" resultid="6234" />
                    <RANKING place="6" resultid="6348" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="13" agemin="12" name="Jahrgang 2010/2011">
                  <RANKINGS>
                    <RANKING place="11" resultid="21" />
                    <RANKING place="18" resultid="150" />
                    <RANKING place="6" resultid="158" />
                    <RANKING place="29" resultid="225" />
                    <RANKING place="2" resultid="612" />
                    <RANKING place="4" resultid="974" />
                    <RANKING place="14" resultid="1915" />
                    <RANKING place="12" resultid="1945" />
                    <RANKING place="28" resultid="1986" />
                    <RANKING place="21" resultid="2033" />
                    <RANKING place="30" resultid="2100" />
                    <RANKING place="31" resultid="2104" />
                    <RANKING place="24" resultid="3759" />
                    <RANKING place="19" resultid="3773" />
                    <RANKING place="16" resultid="3846" />
                    <RANKING place="7" resultid="4390" />
                    <RANKING place="27" resultid="4549" />
                    <RANKING place="15" resultid="4930" />
                    <RANKING place="13" resultid="4933" />
                    <RANKING place="25" resultid="4970" />
                    <RANKING place="20" resultid="5030" />
                    <RANKING place="8" resultid="5151" />
                    <RANKING place="5" resultid="5240" />
                    <RANKING place="9" resultid="5297" />
                    <RANKING place="3" resultid="5393" />
                    <RANKING place="22" resultid="5463" />
                    <RANKING place="1" resultid="5501" />
                    <RANKING place="17" resultid="5557" />
                    <RANKING place="32" resultid="5707" />
                    <RANKING place="23" resultid="5791" />
                    <RANKING place="10" resultid="5801" />
                    <RANKING place="26" resultid="6286" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6" agemax="15" agemin="14" name="Jahrgang 2008/2009">
                  <RANKINGS>
                    <RANKING place="15" resultid="1924" />
                    <RANKING place="14" resultid="3721" />
                    <RANKING place="1" resultid="4582" />
                    <RANKING place="12" resultid="4963" />
                    <RANKING place="13" resultid="4979" />
                    <RANKING place="6" resultid="5274" />
                    <RANKING place="8" resultid="5331" />
                    <RANKING place="2" resultid="5355" />
                    <RANKING place="3" resultid="5433" />
                    <RANKING place="7" resultid="5499" />
                    <RANKING place="4" resultid="5610" />
                    <RANKING place="11" resultid="5652" />
                    <RANKING place="9" resultid="5735" />
                    <RANKING place="10" resultid="5875" />
                    <RANKING place="5" resultid="5915" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8" agemax="17" agemin="16" name="Jahrgang 2006/2007">
                  <RANKINGS>
                    <RANKING place="7" resultid="3745" />
                    <RANKING place="5" resultid="4652" />
                    <RANKING place="3" resultid="4841" />
                    <RANKING place="4" resultid="4961" />
                    <RANKING place="2" resultid="4966" />
                    <RANKING place="6" resultid="4975" />
                    <RANKING place="1" resultid="5488" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="24" number="24" gender="M" round="TIM">
              <SWIMSTYLE stroke="FREE" relaycount="1" distance="200" />
              <HEATS>
                <HEAT heatid="24001" number="1" />
                <HEAT heatid="24002" number="2" />
                <HEAT heatid="24003" number="3" />
                <HEAT heatid="24004" number="4" />
                <HEAT heatid="24005" number="5" />
                <HEAT heatid="24006" number="6" />
                <HEAT heatid="24007" number="7" />
                <HEAT heatid="24008" number="8" />
                <HEAT heatid="24009" number="9" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="10" agemin="10" name="Jahrgang 2013">
                  <RANKINGS>
                    <RANKING place="12" resultid="2130" />
                    <RANKING place="1" resultid="3435" />
                    <RANKING place="5" resultid="4042" />
                    <RANKING place="10" resultid="4250" />
                    <RANKING place="4" resultid="4345" />
                    <RANKING place="3" resultid="4393" />
                    <RANKING place="8" resultid="4762" />
                    <RANKING place="6" resultid="4985" />
                    <RANKING place="9" resultid="5174" />
                    <RANKING place="11" resultid="5539" />
                    <RANKING place="2" resultid="5627" />
                    <RANKING place="7" resultid="5946" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2" agemax="11" agemin="11" name="Jahrgang 2012">
                  <RANKINGS>
                    <RANKING place="1" resultid="126" />
                    <RANKING place="15" resultid="812" />
                    <RANKING place="14" resultid="856" />
                    <RANKING place="9" resultid="915" />
                    <RANKING place="11" resultid="990" />
                    <RANKING place="16" resultid="998" />
                    <RANKING place="7" resultid="2134" />
                    <RANKING place="10" resultid="4068" />
                    <RANKING place="4" resultid="4114" />
                    <RANKING place="5" resultid="4452" />
                    <RANKING place="13" resultid="4720" />
                    <RANKING place="3" resultid="4727" />
                    <RANKING place="12" resultid="4799" />
                    <RANKING place="2" resultid="5171" />
                    <RANKING place="6" resultid="5520" />
                    <RANKING place="8" resultid="5941" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="13" agemin="12" name="Jahrgang 2010/2011">
                  <RANKINGS>
                    <RANKING place="3" resultid="791" />
                    <RANKING place="1" resultid="870" />
                    <RANKING place="24" resultid="1889" />
                    <RANKING place="15" resultid="1984" />
                    <RANKING place="23" resultid="2047" />
                    <RANKING place="21" resultid="3733" />
                    <RANKING place="4" resultid="4469" />
                    <RANKING place="17" resultid="4542" />
                    <RANKING place="16" resultid="4565" />
                    <RANKING place="9" resultid="4594" />
                    <RANKING place="13" resultid="4606" />
                    <RANKING place="19" resultid="4611" />
                    <RANKING place="6" resultid="4630" />
                    <RANKING place="7" resultid="4794" />
                    <RANKING place="11" resultid="4894" />
                    <RANKING place="14" resultid="4989" />
                    <RANKING place="8" resultid="5244" />
                    <RANKING place="18" resultid="5266" />
                    <RANKING place="22" resultid="5513" />
                    <RANKING place="2" resultid="5699" />
                    <RANKING place="5" resultid="5750" />
                    <RANKING place="20" resultid="5898" />
                    <RANKING place="12" resultid="6310" />
                    <RANKING place="10" resultid="6331" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6" agemax="15" agemin="14" name="Jahrgang 2008/2009">
                  <RANKINGS>
                    <RANKING place="8" resultid="3490" />
                    <RANKING place="9" resultid="3769" />
                    <RANKING place="7" resultid="4601" />
                    <RANKING place="5" resultid="4663" />
                    <RANKING place="6" resultid="5069" />
                    <RANKING place="4" resultid="5363" />
                    <RANKING place="3" resultid="5510" />
                    <RANKING place="2" resultid="5902" />
                    <RANKING place="1" resultid="6019" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8" agemax="17" agemin="16" name="Jahrgang 2006/2007">
                  <RANKINGS>
                    <RANKING place="3" resultid="4298" />
                    <RANKING place="1" resultid="5136" />
                    <RANKING place="2" resultid="6307" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="25" number="25" gender="F" round="TIM">
              <SWIMSTYLE stroke="BACK" relaycount="1" distance="50" />
              <HEATS>
                <HEAT heatid="25001" number="1" />
                <HEAT heatid="25002" number="2" />
                <HEAT heatid="25003" number="3" />
                <HEAT heatid="25004" number="4" />
                <HEAT heatid="25005" number="5" />
                <HEAT heatid="25006" number="6" />
                <HEAT heatid="25007" number="7" />
                <HEAT heatid="25008" number="8" />
                <HEAT heatid="25009" number="9" />
                <HEAT heatid="25010" number="10" />
                <HEAT heatid="25011" number="11" />
                <HEAT heatid="25012" number="12" />
                <HEAT heatid="25013" number="13" />
                <HEAT heatid="25014" number="14" />
                <HEAT heatid="25015" number="15" />
                <HEAT heatid="25016" number="16" />
                <HEAT heatid="25017" number="17" />
                <HEAT heatid="25018" number="18" />
                <HEAT heatid="25019" number="19" />
                <HEAT heatid="25020" number="20" />
                <HEAT heatid="25021" number="21" />
                <HEAT heatid="25022" number="22" />
                <HEAT heatid="25023" number="23" />
                <HEAT heatid="25024" number="24" />
                <HEAT heatid="25025" number="25" />
                <HEAT heatid="25026" number="26" />
                <HEAT heatid="25027" number="27" />
                <HEAT heatid="25028" number="28" />
                <HEAT heatid="25029" number="29" />
                <HEAT heatid="25030" number="30" />
                <HEAT heatid="25031" number="31" />
                <HEAT heatid="25032" number="32" />
                <HEAT heatid="25033" number="33" />
                <HEAT heatid="25034" number="34" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="10" agemax="8" agemin="8" name="Jahrgang 2015">
                  <RANKINGS>
                    <RANKING place="9" resultid="199" />
                    <RANKING place="10" resultid="222" />
                    <RANKING place="48" resultid="866" />
                    <RANKING place="12" resultid="877" />
                    <RANKING place="42" resultid="901" />
                    <RANKING place="41" resultid="905" />
                    <RANKING place="35" resultid="1005" />
                    <RANKING place="51" resultid="1901" />
                    <RANKING place="52" resultid="1926" />
                    <RANKING place="16" resultid="1973" />
                    <RANKING place="21" resultid="1979" />
                    <RANKING place="6" resultid="2075" />
                    <RANKING place="5" resultid="3448" />
                    <RANKING place="22" resultid="3831" />
                    <RANKING place="49" resultid="4057" />
                    <RANKING place="25" resultid="4090" />
                    <RANKING place="20" resultid="4155" />
                    <RANKING place="8" resultid="4203" />
                    <RANKING place="23" resultid="4220" />
                    <RANKING place="11" resultid="4224" />
                    <RANKING place="28" resultid="4253" />
                    <RANKING place="4" resultid="4338" />
                    <RANKING place="44" resultid="4352" />
                    <RANKING place="14" resultid="4386" />
                    <RANKING place="26" resultid="4449" />
                    <RANKING place="33" resultid="4472" />
                    <RANKING place="13" resultid="4490" />
                    <RANKING place="24" resultid="4527" />
                    <RANKING place="46" resultid="4587" />
                    <RANKING place="45" resultid="4755" />
                    <RANKING place="50" resultid="4938" />
                    <RANKING place="29" resultid="5007" />
                    <RANKING place="43" resultid="5042" />
                    <RANKING place="34" resultid="5056" />
                    <RANKING place="35" resultid="5074" />
                    <RANKING place="17" resultid="5092" />
                    <RANKING place="7" resultid="5119" />
                    <RANKING place="47" resultid="5124" />
                    <RANKING place="2" resultid="5128" />
                    <RANKING place="15" resultid="5202" />
                    <RANKING place="19" resultid="5226" />
                    <RANKING place="38" resultid="5857" />
                    <RANKING place="1" resultid="5967" />
                    <RANKING place="18" resultid="5982" />
                    <RANKING place="26" resultid="6076" />
                    <RANKING place="31" resultid="6091" />
                    <RANKING place="32" resultid="6112" />
                    <RANKING place="39" resultid="6130" />
                    <RANKING place="40" resultid="6134" />
                    <RANKING place="29" resultid="6174" />
                    <RANKING place="37" resultid="6230" />
                    <RANKING place="3" resultid="6297" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9" agemax="9" agemin="9" name="Jahrgang 2014">
                  <RANKINGS>
                    <RANKING place="56" resultid="229" />
                    <RANKING place="60" resultid="837" />
                    <RANKING place="43" resultid="910" />
                    <RANKING place="25" resultid="935" />
                    <RANKING place="2" resultid="965" />
                    <RANKING place="21" resultid="1636" />
                    <RANKING place="3" resultid="1641" />
                    <RANKING place="28" resultid="1657" />
                    <RANKING place="19" resultid="1661" />
                    <RANKING place="31" resultid="1907" />
                    <RANKING place="58" resultid="1941" />
                    <RANKING place="27" resultid="2015" />
                    <RANKING place="32" resultid="2095" />
                    <RANKING place="24" resultid="3451" />
                    <RANKING place="12" resultid="3479" />
                    <RANKING place="59" resultid="3718" />
                    <RANKING place="46" resultid="4084" />
                    <RANKING place="54" resultid="4094" />
                    <RANKING place="42" resultid="4140" />
                    <RANKING place="48" resultid="4275" />
                    <RANKING place="1" resultid="4279" />
                    <RANKING place="47" resultid="4306" />
                    <RANKING place="40" resultid="4310" />
                    <RANKING place="38" resultid="4328" />
                    <RANKING place="15" resultid="4333" />
                    <RANKING place="17" resultid="4363" />
                    <RANKING place="37" resultid="4372" />
                    <RANKING place="8" resultid="4381" />
                    <RANKING place="13" resultid="4410" />
                    <RANKING place="29" resultid="4433" />
                    <RANKING place="18" resultid="4461" />
                    <RANKING place="61" resultid="4645" />
                    <RANKING place="35" resultid="4766" />
                    <RANKING place="55" resultid="5020" />
                    <RANKING place="22" resultid="5078" />
                    <RANKING place="36" resultid="5102" />
                    <RANKING place="50" resultid="5113" />
                    <RANKING place="14" resultid="5214" />
                    <RANKING place="44" resultid="5292" />
                    <RANKING place="8" resultid="5377" />
                    <RANKING place="39" resultid="5398" />
                    <RANKING place="52" resultid="5448" />
                    <RANKING place="20" resultid="5483" />
                    <RANKING place="57" resultid="5508" />
                    <RANKING place="51" resultid="5533" />
                    <RANKING place="33" resultid="5553" />
                    <RANKING place="41" resultid="5560" />
                    <RANKING place="30" resultid="5596" />
                    <RANKING place="23" resultid="5632" />
                    <RANKING place="7" resultid="5678" />
                    <RANKING place="45" resultid="5756" />
                    <RANKING place="49" resultid="5863" />
                    <RANKING place="4" resultid="5866" />
                    <RANKING place="53" resultid="5869" />
                    <RANKING place="5" resultid="5907" />
                    <RANKING place="34" resultid="6056" />
                    <RANKING place="6" resultid="6060" />
                    <RANKING place="10" resultid="6151" />
                    <RANKING place="11" resultid="6194" />
                    <RANKING place="16" resultid="6214" />
                    <RANKING place="25" resultid="6290" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1" agemax="10" agemin="10" name="Jahrgang 2013">
                  <RANKINGS>
                    <RANKING place="1" resultid="11" />
                    <RANKING place="10" resultid="213" />
                    <RANKING place="12" resultid="247" />
                    <RANKING place="13" resultid="474" />
                    <RANKING place="17" resultid="762" />
                    <RANKING place="4" resultid="765" />
                    <RANKING place="2" resultid="798" />
                    <RANKING place="11" resultid="886" />
                    <RANKING place="28" resultid="948" />
                    <RANKING place="8" resultid="1918" />
                    <RANKING place="31" resultid="1964" />
                    <RANKING place="26" resultid="1997" />
                    <RANKING place="19" resultid="3492" />
                    <RANKING place="25" resultid="3728" />
                    <RANKING place="16" resultid="4358" />
                    <RANKING place="9" resultid="4445" />
                    <RANKING place="15" resultid="4456" />
                    <RANKING place="13" resultid="4474" />
                    <RANKING place="23" resultid="4637" />
                    <RANKING place="20" resultid="4750" />
                    <RANKING place="22" resultid="5097" />
                    <RANKING place="5" resultid="5143" />
                    <RANKING place="18" resultid="5193" />
                    <RANKING place="6" resultid="5223" />
                    <RANKING place="24" resultid="5249" />
                    <RANKING place="3" resultid="5443" />
                    <RANKING place="30" resultid="5772" />
                    <RANKING place="29" resultid="5782" />
                    <RANKING place="21" resultid="6052" />
                    <RANKING place="7" resultid="6108" />
                    <RANKING place="27" resultid="6325" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2" agemax="11" agemin="11" name="Jahrgang 2012">
                  <RANKINGS>
                    <RANKING place="8" resultid="19" />
                    <RANKING place="18" resultid="182" />
                    <RANKING place="15" resultid="806" />
                    <RANKING place="4" resultid="956" />
                    <RANKING place="9" resultid="1596" />
                    <RANKING place="13" resultid="1607" />
                    <RANKING place="25" resultid="1891" />
                    <RANKING place="21" resultid="1949" />
                    <RANKING place="5" resultid="1991" />
                    <RANKING place="28" resultid="3811" />
                    <RANKING place="30" resultid="4479" />
                    <RANKING place="14" resultid="4508" />
                    <RANKING place="35" resultid="4562" />
                    <RANKING place="10" resultid="4741" />
                    <RANKING place="19" resultid="4815" />
                    <RANKING place="7" resultid="4914" />
                    <RANKING place="24" resultid="4921" />
                    <RANKING place="22" resultid="5037" />
                    <RANKING place="29" resultid="5109" />
                    <RANKING place="11" resultid="5233" />
                    <RANKING place="1" resultid="5344" />
                    <RANKING place="23" resultid="5494" />
                    <RANKING place="33" resultid="5621" />
                    <RANKING place="16" resultid="5646" />
                    <RANKING place="26" resultid="5673" />
                    <RANKING place="2" resultid="5714" />
                    <RANKING place="17" resultid="5722" />
                    <RANKING place="32" resultid="5796" />
                    <RANKING place="36" resultid="5819" />
                    <RANKING place="11" resultid="5845" />
                    <RANKING place="34" resultid="5860" />
                    <RANKING place="20" resultid="5975" />
                    <RANKING place="3" resultid="6038" />
                    <RANKING place="27" resultid="6304" />
                    <RANKING place="6" resultid="6335" />
                    <RANKING place="31" resultid="6341" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="13" agemin="12" name="Jahrgang 2010/2011">
                  <RANKINGS>
                    <RANKING place="10" resultid="22" />
                    <RANKING place="1" resultid="134" />
                    <RANKING place="7" resultid="174" />
                    <RANKING place="30" resultid="226" />
                    <RANKING place="3" resultid="973" />
                    <RANKING place="13" resultid="2060" />
                    <RANKING place="29" resultid="2099" />
                    <RANKING place="18" resultid="2103" />
                    <RANKING place="8" resultid="2138" />
                    <RANKING place="37" resultid="3740" />
                    <RANKING place="39" resultid="3753" />
                    <RANKING place="40" resultid="3779" />
                    <RANKING place="35" resultid="4302" />
                    <RANKING place="23" resultid="4391" />
                    <RANKING place="9" resultid="4443" />
                    <RANKING place="21" resultid="4550" />
                    <RANKING place="31" resultid="4560" />
                    <RANKING place="15" resultid="4698" />
                    <RANKING place="17" resultid="4847" />
                    <RANKING place="12" resultid="4868" />
                    <RANKING place="22" resultid="4882" />
                    <RANKING place="26" resultid="4931" />
                    <RANKING place="14" resultid="4934" />
                    <RANKING place="16" resultid="4971" />
                    <RANKING place="36" resultid="5003" />
                    <RANKING place="25" resultid="5031" />
                    <RANKING place="20" resultid="5087" />
                    <RANKING place="19" resultid="5149" />
                    <RANKING place="6" resultid="5210" />
                    <RANKING place="4" resultid="5241" />
                    <RANKING place="11" resultid="5298" />
                    <RANKING place="33" resultid="5371" />
                    <RANKING place="2" resultid="5394" />
                    <RANKING place="5" resultid="5405" />
                    <RANKING place="38" resultid="5505" />
                    <RANKING place="34" resultid="5550" />
                    <RANKING place="27" resultid="5607" />
                    <RANKING place="32" resultid="5708" />
                    <RANKING place="28" resultid="5763" />
                    <RANKING place="24" resultid="6287" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6" agemax="15" agemin="14" name="Jahrgang 2008/2009">
                  <RANKINGS>
                    <RANKING place="20" resultid="1923" />
                    <RANKING place="1" resultid="2011" />
                    <RANKING place="16" resultid="3460" />
                    <RANKING place="6" resultid="4291" />
                    <RANKING place="3" resultid="4583" />
                    <RANKING place="15" resultid="4745" />
                    <RANKING place="11" resultid="4888" />
                    <RANKING place="7" resultid="4944" />
                    <RANKING place="13" resultid="4964" />
                    <RANKING place="14" resultid="4980" />
                    <RANKING place="4" resultid="4996" />
                    <RANKING place="18" resultid="5275" />
                    <RANKING place="17" resultid="5295" />
                    <RANKING place="9" resultid="5332" />
                    <RANKING place="5" resultid="5356" />
                    <RANKING place="19" resultid="5666" />
                    <RANKING place="10" resultid="5736" />
                    <RANKING place="12" resultid="5922" />
                    <RANKING place="2" resultid="6140" />
                    <RANKING place="8" resultid="6159" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8" agemax="17" agemin="16" name="Jahrgang 2006/2007">
                  <RANKINGS>
                    <RANKING place="2" resultid="3726" />
                    <RANKING place="5" resultid="3809" />
                    <RANKING place="3" resultid="4731" />
                    <RANKING place="1" resultid="4967" />
                    <RANKING place="4" resultid="4976" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="26" number="26" gender="M" round="TIM">
              <SWIMSTYLE stroke="BACK" relaycount="1" distance="50" />
              <HEATS>
                <HEAT heatid="26001" number="1" />
                <HEAT heatid="26002" number="2" />
                <HEAT heatid="26003" number="3" />
                <HEAT heatid="26004" number="4" />
                <HEAT heatid="26005" number="5" />
                <HEAT heatid="26006" number="6" />
                <HEAT heatid="26007" number="7" />
                <HEAT heatid="26008" number="8" />
                <HEAT heatid="26009" number="9" />
                <HEAT heatid="26010" number="10" />
                <HEAT heatid="26011" number="11" />
                <HEAT heatid="26012" number="12" />
                <HEAT heatid="26013" number="13" />
                <HEAT heatid="26014" number="14" />
                <HEAT heatid="26015" number="15" />
                <HEAT heatid="26016" number="16" />
                <HEAT heatid="26017" number="17" />
                <HEAT heatid="26018" number="18" />
                <HEAT heatid="26019" number="19" />
                <HEAT heatid="26020" number="20" />
                <HEAT heatid="26021" number="21" />
                <HEAT heatid="26022" number="22" />
                <HEAT heatid="26023" number="23" />
                <HEAT heatid="26024" number="24" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="10" agemax="8" agemin="8" name="Jahrgang 2015">
                  <RANKINGS>
                    <RANKING place="33" resultid="195" />
                    <RANKING place="19" resultid="206" />
                    <RANKING place="30" resultid="833" />
                    <RANKING place="32" resultid="930" />
                    <RANKING place="16" resultid="938" />
                    <RANKING place="7" resultid="968" />
                    <RANKING place="20" resultid="1884" />
                    <RANKING place="23" resultid="1897" />
                    <RANKING place="6" resultid="2028" />
                    <RANKING place="21" resultid="2066" />
                    <RANKING place="24" resultid="4081" />
                    <RANKING place="22" resultid="4165" />
                    <RANKING place="5" resultid="4186" />
                    <RANKING place="1" resultid="4378" />
                    <RANKING place="8" resultid="4494" />
                    <RANKING place="9" resultid="4519" />
                    <RANKING place="4" resultid="4524" />
                    <RANKING place="14" resultid="4681" />
                    <RANKING place="11" resultid="4714" />
                    <RANKING place="26" resultid="4790" />
                    <RANKING place="3" resultid="5017" />
                    <RANKING place="2" resultid="5655" />
                    <RANKING place="29" resultid="5971" />
                    <RANKING place="31" resultid="5985" />
                    <RANKING place="18" resultid="5989" />
                    <RANKING place="25" resultid="5993" />
                    <RANKING place="12" resultid="6016" />
                    <RANKING place="28" resultid="6068" />
                    <RANKING place="13" resultid="6105" />
                    <RANKING place="15" resultid="6164" />
                    <RANKING place="17" resultid="6205" />
                    <RANKING place="10" resultid="6208" />
                    <RANKING place="27" resultid="6227" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9" agemax="9" agemin="9" name="Jahrgang 2014">
                  <RANKINGS>
                    <RANKING place="25" resultid="238" />
                    <RANKING place="29" resultid="479" />
                    <RANKING place="5" resultid="882" />
                    <RANKING place="36" resultid="926" />
                    <RANKING place="26" resultid="981" />
                    <RANKING place="37" resultid="986" />
                    <RANKING place="33" resultid="1009" />
                    <RANKING place="3" resultid="1019" />
                    <RANKING place="18" resultid="1603" />
                    <RANKING place="14" resultid="1969" />
                    <RANKING place="11" resultid="2001" />
                    <RANKING place="30" resultid="2050" />
                    <RANKING place="2" resultid="2056" />
                    <RANKING place="9" resultid="4034" />
                    <RANKING place="10" resultid="4047" />
                    <RANKING place="4" resultid="4193" />
                    <RANKING place="13" resultid="4198" />
                    <RANKING place="8" resultid="4207" />
                    <RANKING place="1" resultid="4231" />
                    <RANKING place="24" resultid="4238" />
                    <RANKING place="31" resultid="4655" />
                    <RANKING place="16" resultid="4771" />
                    <RANKING place="22" resultid="5050" />
                    <RANKING place="17" resultid="5185" />
                    <RANKING place="27" resultid="5197" />
                    <RANKING place="19" resultid="5408" />
                    <RANKING place="20" resultid="5469" />
                    <RANKING place="7" resultid="5601" />
                    <RANKING place="15" resultid="5695" />
                    <RANKING place="6" resultid="5730" />
                    <RANKING place="32" resultid="6155" />
                    <RANKING place="12" resultid="6218" />
                    <RANKING place="34" resultid="6256" />
                    <RANKING place="23" resultid="6280" />
                    <RANKING place="28" resultid="6343" />
                    <RANKING place="35" resultid="6355" />
                    <RANKING place="21" resultid="6358" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1" agemax="10" agemin="10" name="Jahrgang 2013">
                  <RANKINGS>
                    <RANKING place="11" resultid="759" />
                    <RANKING place="1" resultid="943" />
                    <RANKING place="18" resultid="2035" />
                    <RANKING place="23" resultid="3496" />
                    <RANKING place="21" resultid="3736" />
                    <RANKING place="12" resultid="4053" />
                    <RANKING place="9" resultid="4101" />
                    <RANKING place="10" resultid="4178" />
                    <RANKING place="13" resultid="4422" />
                    <RANKING place="5" resultid="4498" />
                    <RANKING place="15" resultid="4763" />
                    <RANKING place="16" resultid="4779" />
                    <RANKING place="8" resultid="4986" />
                    <RANKING place="17" resultid="5065" />
                    <RANKING place="22" resultid="5544" />
                    <RANKING place="14" resultid="5589" />
                    <RANKING place="4" resultid="5838" />
                    <RANKING place="3" resultid="5891" />
                    <RANKING place="2" resultid="5954" />
                    <RANKING place="7" resultid="6200" />
                    <RANKING place="6" resultid="6263" />
                    <RANKING place="19" resultid="6268" />
                    <RANKING place="20" resultid="6314" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2" agemax="11" agemin="11" name="Jahrgang 2012">
                  <RANKINGS>
                    <RANKING place="1" resultid="190" />
                    <RANKING place="24" resultid="203" />
                    <RANKING place="13" resultid="783" />
                    <RANKING place="9" resultid="819" />
                    <RANKING place="15" resultid="914" />
                    <RANKING place="6" resultid="3456" />
                    <RANKING place="14" resultid="4069" />
                    <RANKING place="18" resultid="4271" />
                    <RANKING place="16" resultid="4349" />
                    <RANKING place="11" resultid="4418" />
                    <RANKING place="5" resultid="4728" />
                    <RANKING place="12" resultid="4828" />
                    <RANKING place="3" resultid="5172" />
                    <RANKING place="21" resultid="5310" />
                    <RANKING place="4" resultid="5521" />
                    <RANKING place="8" resultid="5528" />
                    <RANKING place="20" resultid="5570" />
                    <RANKING place="7" resultid="5690" />
                    <RANKING place="17" resultid="5806" />
                    <RANKING place="25" resultid="5812" />
                    <RANKING place="19" resultid="5853" />
                    <RANKING place="10" resultid="5942" />
                    <RANKING place="2" resultid="6185" />
                    <RANKING place="23" resultid="6253" />
                    <RANKING place="22" resultid="6272" />
                    <RANKING place="26" resultid="6301" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="13" agemin="12" name="Jahrgang 2010/2011">
                  <RANKINGS>
                    <RANKING place="3" resultid="118" />
                    <RANKING place="5" resultid="142" />
                    <RANKING place="2" resultid="769" />
                    <RANKING place="1" resultid="809" />
                    <RANKING place="31" resultid="1888" />
                    <RANKING place="11" resultid="1930" />
                    <RANKING place="20" resultid="2046" />
                    <RANKING place="18" resultid="2089" />
                    <RANKING place="6" resultid="3441" />
                    <RANKING place="33" resultid="3847" />
                    <RANKING place="9" resultid="4288" />
                    <RANKING place="19" resultid="4543" />
                    <RANKING place="27" resultid="4555" />
                    <RANKING place="30" resultid="4566" />
                    <RANKING place="21" resultid="4572" />
                    <RANKING place="23" resultid="4607" />
                    <RANKING place="25" resultid="4612" />
                    <RANKING place="28" resultid="4642" />
                    <RANKING place="14" resultid="4895" />
                    <RANKING place="22" resultid="4902" />
                    <RANKING place="15" resultid="4990" />
                    <RANKING place="8" resultid="5245" />
                    <RANKING place="24" resultid="5267" />
                    <RANKING place="7" resultid="5427" />
                    <RANKING place="29" resultid="5514" />
                    <RANKING place="32" resultid="5593" />
                    <RANKING place="13" resultid="5662" />
                    <RANKING place="4" resultid="5751" />
                    <RANKING place="10" resultid="5884" />
                    <RANKING place="16" resultid="5899" />
                    <RANKING place="12" resultid="6167" />
                    <RANKING place="26" resultid="6311" />
                    <RANKING place="17" resultid="6332" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6" agemax="15" agemin="14" name="Jahrgang 2008/2009">
                  <RANKINGS>
                    <RANKING place="9" resultid="3489" />
                    <RANKING place="6" resultid="3774" />
                    <RANKING place="11" resultid="3834" />
                    <RANKING place="12" resultid="4264" />
                    <RANKING place="2" resultid="4318" />
                    <RANKING place="8" resultid="4602" />
                    <RANKING place="13" resultid="4808" />
                    <RANKING place="14" resultid="4822" />
                    <RANKING place="3" resultid="4854" />
                    <RANKING place="5" resultid="4908" />
                    <RANKING place="7" resultid="5070" />
                    <RANKING place="4" resultid="5387" />
                    <RANKING place="1" resultid="6000" />
                    <RANKING place="10" resultid="6083" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8" agemax="17" agemin="16" name="Jahrgang 2006/2007">
                  <RANKINGS>
                    <RANKING place="2" resultid="3464" />
                    <RANKING place="4" resultid="3483" />
                    <RANKING place="3" resultid="3784" />
                    <RANKING place="6" resultid="4835" />
                    <RANKING place="1" resultid="5316" />
                    <RANKING place="7" resultid="5373" />
                    <RANKING place="5" resultid="6308" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="27" number="27" gender="F" round="TIM">
              <SWIMSTYLE stroke="BREAST" name="50 Brustbeinbewegung Frauen" technique="KICK" relaycount="1" distance="50" />
              <HEATS>
                <HEAT heatid="27000" number="0" />
                <HEAT heatid="27001" number="1" />
                <HEAT heatid="27002" number="2" />
                <HEAT heatid="27003" number="3" />
                <HEAT heatid="27004" number="4" />
                <HEAT heatid="27005" number="5" />
                <HEAT heatid="27006" number="6" />
                <HEAT heatid="27007" number="7" />
                <HEAT heatid="27008" number="8" />
                <HEAT heatid="27009" number="9" />
                <HEAT heatid="27010" number="10" />
                <HEAT heatid="27011" number="11" />
                <HEAT heatid="27012" number="12" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="10" agemax="8" agemin="8" name="Jahrgang 2015">
                  <RANKINGS>
                    <RANKING place="19" resultid="900" />
                    <RANKING place="20" resultid="904" />
                    <RANKING place="15" resultid="1004" />
                    <RANKING place="14" resultid="1900" />
                    <RANKING place="24" resultid="1925" />
                    <RANKING place="26" resultid="1978" />
                    <RANKING place="11" resultid="2074" />
                    <RANKING place="2" resultid="3447" />
                    <RANKING place="7" resultid="3830" />
                    <RANKING place="25" resultid="4058" />
                    <RANKING place="12" resultid="4091" />
                    <RANKING place="18" resultid="4229" />
                    <RANKING place="16" resultid="4254" />
                    <RANKING place="4" resultid="4342" />
                    <RANKING place="9" resultid="4426" />
                    <RANKING place="6" resultid="4450" />
                    <RANKING place="13" resultid="4487" />
                    <RANKING place="3" resultid="4491" />
                    <RANKING place="23" resultid="4528" />
                    <RANKING place="8" resultid="4588" />
                    <RANKING place="30" resultid="4939" />
                    <RANKING place="27" resultid="5008" />
                    <RANKING place="29" resultid="5057" />
                    <RANKING place="28" resultid="5075" />
                    <RANKING place="22" resultid="5120" />
                    <RANKING place="10" resultid="5129" />
                    <RANKING place="5" resultid="5203" />
                    <RANKING place="17" resultid="6009" />
                    <RANKING place="21" resultid="6231" />
                    <RANKING place="1" resultid="6298" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9" agemax="9" agemin="9" name="Jahrgang 2014">
                  <RANKINGS>
                    <RANKING place="1" resultid="802" />
                    <RANKING place="12" resultid="921" />
                    <RANKING place="6" resultid="934" />
                    <RANKING place="22" resultid="1940" />
                    <RANKING place="15" resultid="2069" />
                    <RANKING place="4" resultid="3478" />
                    <RANKING place="20" resultid="3717" />
                    <RANKING place="23" resultid="4150" />
                    <RANKING place="2" resultid="4280" />
                    <RANKING place="5" resultid="4311" />
                    <RANKING place="14" resultid="4364" />
                    <RANKING place="8" resultid="4411" />
                    <RANKING place="19" resultid="5026" />
                    <RANKING place="21" resultid="5045" />
                    <RANKING place="11" resultid="5114" />
                    <RANKING place="9" resultid="5378" />
                    <RANKING place="7" resultid="5449" />
                    <RANKING place="13" resultid="5484" />
                    <RANKING place="24" resultid="5509" />
                    <RANKING place="18" resultid="5534" />
                    <RANKING place="3" resultid="5633" />
                    <RANKING place="10" resultid="5757" />
                    <RANKING place="25" resultid="5870" />
                    <RANKING place="17" resultid="6145" />
                    <RANKING place="16" resultid="6195" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1" agemax="10" agemin="10" name="Jahrgang 2013">
                  <RANKINGS>
                    <RANKING place="3" resultid="780" />
                    <RANKING place="7" resultid="1996" />
                    <RANKING place="6" resultid="3825" />
                    <RANKING place="10" resultid="4130" />
                    <RANKING place="12" resultid="4162" />
                    <RANKING place="5" resultid="4355" />
                    <RANKING place="2" resultid="4457" />
                    <RANKING place="11" resultid="4619" />
                    <RANKING place="4" resultid="5098" />
                    <RANKING place="8" resultid="5466" />
                    <RANKING place="9" resultid="5783" />
                    <RANKING place="1" resultid="5832" />
                    <RANKING place="13" resultid="5928" />
                    <RANKING place="14" resultid="6046" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2" agemax="11" agemin="11" name="Jahrgang 2012">
                  <RANKINGS>
                    <RANKING place="10" resultid="1645" />
                    <RANKING place="14" resultid="4563" />
                    <RANKING place="5" resultid="4816" />
                    <RANKING place="6" resultid="4875" />
                    <RANKING place="4" resultid="5038" />
                    <RANKING place="9" resultid="5674" />
                    <RANKING place="8" resultid="5723" />
                    <RANKING place="13" resultid="5797" />
                    <RANKING place="7" resultid="5861" />
                    <RANKING place="2" resultid="6027" />
                    <RANKING place="12" resultid="6180" />
                    <RANKING place="3" resultid="6235" />
                    <RANKING place="11" resultid="6305" />
                    <RANKING place="15" resultid="6336" />
                    <RANKING place="1" resultid="6365" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="28" number="28" gender="M" round="TIM">
              <SWIMSTYLE stroke="BREAST" name="50 Brustbeinbewegung Männer" technique="KICK" relaycount="1" distance="50" />
              <HEATS>
                <HEAT heatid="28001" number="1" />
                <HEAT heatid="28002" number="2" />
                <HEAT heatid="28003" number="3" />
                <HEAT heatid="28004" number="4" />
                <HEAT heatid="28005" number="5" />
                <HEAT heatid="28006" number="6" />
                <HEAT heatid="28007" number="7" />
                <HEAT heatid="28008" number="8" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="10" agemax="8" agemin="8" name="Jahrgang 2015">
                  <RANKINGS>
                    <RANKING place="6" resultid="862" />
                    <RANKING place="15" resultid="929" />
                    <RANKING place="8" resultid="1896" />
                    <RANKING place="13" resultid="2027" />
                    <RANKING place="2" resultid="3842" />
                    <RANKING place="9" resultid="4082" />
                    <RANKING place="1" resultid="4398" />
                    <RANKING place="3" resultid="4495" />
                    <RANKING place="7" resultid="4520" />
                    <RANKING place="4" resultid="4924" />
                    <RANKING place="5" resultid="5656" />
                    <RANKING place="10" resultid="5986" />
                    <RANKING place="12" resultid="6069" />
                    <RANKING place="11" resultid="6072" />
                    <RANKING place="14" resultid="6123" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9" agemax="9" agemin="9" name="Jahrgang 2014">
                  <RANKINGS>
                    <RANKING place="9" resultid="480" />
                    <RANKING place="9" resultid="925" />
                    <RANKING place="16" resultid="980" />
                    <RANKING place="17" resultid="985" />
                    <RANKING place="19" resultid="1008" />
                    <RANKING place="2" resultid="1018" />
                    <RANKING place="13" resultid="1620" />
                    <RANKING place="15" resultid="2019" />
                    <RANKING place="4" resultid="4191" />
                    <RANKING place="6" resultid="4199" />
                    <RANKING place="1" resultid="4211" />
                    <RANKING place="12" resultid="4534" />
                    <RANKING place="18" resultid="4656" />
                    <RANKING place="5" resultid="5409" />
                    <RANKING place="7" resultid="5696" />
                    <RANKING place="3" resultid="5731" />
                    <RANKING place="20" resultid="5959" />
                    <RANKING place="11" resultid="5997" />
                    <RANKING place="8" resultid="6243" />
                    <RANKING place="14" resultid="6344" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1" agemax="10" agemin="10" name="Jahrgang 2013">
                  <RANKINGS>
                    <RANKING place="3" resultid="849" />
                    <RANKING place="5" resultid="1622" />
                    <RANKING place="4" resultid="1629" />
                    <RANKING place="8" resultid="3495" />
                    <RANKING place="10" resultid="3838" />
                    <RANKING place="2" resultid="4367" />
                    <RANKING place="6" resultid="4499" />
                    <RANKING place="9" resultid="5066" />
                    <RANKING place="11" resultid="5545" />
                    <RANKING place="1" resultid="5590" />
                    <RANKING place="7" resultid="6201" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2" agemax="11" agemin="11" name="Jahrgang 2012">
                  <RANKINGS>
                    <RANKING place="4" resultid="166" />
                    <RANKING place="2" resultid="2006" />
                    <RANKING place="10" resultid="3747" />
                    <RANKING place="8" resultid="3787" />
                    <RANKING place="3" resultid="4243" />
                    <RANKING place="1" resultid="4401" />
                    <RANKING place="7" resultid="4482" />
                    <RANKING place="6" resultid="4829" />
                    <RANKING place="9" resultid="5813" />
                    <RANKING place="5" resultid="6011" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="29" number="29" gender="F" round="TIM">
              <SWIMSTYLE stroke="FREE" relaycount="1" distance="50" />
              <HEATS>
                <HEAT heatid="29001" number="1" />
                <HEAT heatid="29002" number="2" />
                <HEAT heatid="29003" number="3" />
                <HEAT heatid="29004" number="4" />
                <HEAT heatid="29005" number="5" />
                <HEAT heatid="29006" number="6" />
                <HEAT heatid="29007" number="7" />
                <HEAT heatid="29008" number="8" />
                <HEAT heatid="29009" number="9" />
                <HEAT heatid="29010" number="10" />
                <HEAT heatid="29011" number="11" />
                <HEAT heatid="29012" number="12" />
                <HEAT heatid="29013" number="13" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="10" agemax="8" agemin="8" name="Jahrgang 2015">
                  <RANKINGS>
                    <RANKING place="35" resultid="865" />
                    <RANKING place="11" resultid="876" />
                    <RANKING place="36" resultid="899" />
                    <RANKING place="20" resultid="903" />
                    <RANKING place="33" resultid="1003" />
                    <RANKING place="15" resultid="1972" />
                    <RANKING place="25" resultid="1977" />
                    <RANKING place="12" resultid="2073" />
                    <RANKING place="5" resultid="3446" />
                    <RANKING place="32" resultid="3829" />
                    <RANKING place="34" resultid="4092" />
                    <RANKING place="14" resultid="4156" />
                    <RANKING place="31" resultid="4204" />
                    <RANKING place="28" resultid="4221" />
                    <RANKING place="10" resultid="4225" />
                    <RANKING place="21" resultid="4255" />
                    <RANKING place="2" resultid="4339" />
                    <RANKING place="8" resultid="4343" />
                    <RANKING place="3" resultid="4387" />
                    <RANKING place="26" resultid="4416" />
                    <RANKING place="18" resultid="4427" />
                    <RANKING place="23" resultid="4488" />
                    <RANKING place="9" resultid="4492" />
                    <RANKING place="16" resultid="4529" />
                    <RANKING place="27" resultid="5009" />
                    <RANKING place="19" resultid="5043" />
                    <RANKING place="24" resultid="5076" />
                    <RANKING place="7" resultid="5093" />
                    <RANKING place="6" resultid="5121" />
                    <RANKING place="30" resultid="5125" />
                    <RANKING place="1" resultid="5130" />
                    <RANKING place="13" resultid="5204" />
                    <RANKING place="22" resultid="5227" />
                    <RANKING place="4" resultid="5968" />
                    <RANKING place="17" resultid="5983" />
                    <RANKING place="29" resultid="6113" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9" agemax="9" agemin="9" name="Jahrgang 2014">
                  <RANKINGS>
                    <RANKING place="9" resultid="801" />
                    <RANKING place="58" resultid="836" />
                    <RANKING place="44" resultid="909" />
                    <RANKING place="25" resultid="920" />
                    <RANKING place="52" resultid="933" />
                    <RANKING place="2" resultid="964" />
                    <RANKING place="13" resultid="1635" />
                    <RANKING place="3" resultid="1640" />
                    <RANKING place="8" resultid="1656" />
                    <RANKING place="21" resultid="1660" />
                    <RANKING place="26" resultid="1906" />
                    <RANKING place="60" resultid="1939" />
                    <RANKING place="49" resultid="2014" />
                    <RANKING place="56" resultid="2068" />
                    <RANKING place="51" resultid="2094" />
                    <RANKING place="19" resultid="3450" />
                    <RANKING place="39" resultid="4085" />
                    <RANKING place="47" resultid="4095" />
                    <RANKING place="6" resultid="4122" />
                    <RANKING place="37" resultid="4141" />
                    <RANKING place="48" resultid="4151" />
                    <RANKING place="18" resultid="4276" />
                    <RANKING place="1" resultid="4281" />
                    <RANKING place="38" resultid="4307" />
                    <RANKING place="43" resultid="4312" />
                    <RANKING place="12" resultid="4329" />
                    <RANKING place="33" resultid="4334" />
                    <RANKING place="16" resultid="4373" />
                    <RANKING place="7" resultid="4382" />
                    <RANKING place="14" resultid="4434" />
                    <RANKING place="29" resultid="4462" />
                    <RANKING place="61" resultid="4646" />
                    <RANKING place="22" resultid="4767" />
                    <RANKING place="50" resultid="5022" />
                    <RANKING place="40" resultid="5027" />
                    <RANKING place="32" resultid="5046" />
                    <RANKING place="11" resultid="5079" />
                    <RANKING place="27" resultid="5103" />
                    <RANKING place="42" resultid="5115" />
                    <RANKING place="15" resultid="5215" />
                    <RANKING place="34" resultid="5293" />
                    <RANKING place="16" resultid="5379" />
                    <RANKING place="5" resultid="5383" />
                    <RANKING place="46" resultid="5399" />
                    <RANKING place="54" resultid="5450" />
                    <RANKING place="41" resultid="5535" />
                    <RANKING place="31" resultid="5554" />
                    <RANKING place="28" resultid="5561" />
                    <RANKING place="45" resultid="5597" />
                    <RANKING place="35" resultid="5634" />
                    <RANKING place="20" resultid="5679" />
                    <RANKING place="4" resultid="5867" />
                    <RANKING place="57" resultid="5871" />
                    <RANKING place="30" resultid="5908" />
                    <RANKING place="53" resultid="6057" />
                    <RANKING place="36" resultid="6061" />
                    <RANKING place="55" resultid="6086" />
                    <RANKING place="24" resultid="6146" />
                    <RANKING place="59" resultid="6147" />
                    <RANKING place="23" resultid="6152" />
                    <RANKING place="10" resultid="6215" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="30" number="30" gender="M" round="TIM">
              <SWIMSTYLE stroke="FREE" relaycount="1" distance="50" />
              <HEATS>
                <HEAT heatid="30001" number="1" />
                <HEAT heatid="30002" number="2" />
                <HEAT heatid="30003" number="3" />
                <HEAT heatid="30004" number="4" />
                <HEAT heatid="30005" number="5" />
                <HEAT heatid="30006" number="6" />
                <HEAT heatid="30007" number="7" />
                <HEAT heatid="30008" number="8" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="10" agemax="8" agemin="8" name="Jahrgang 2015">
                  <RANKINGS>
                    <RANKING place="23" resultid="832" />
                    <RANKING place="19" resultid="861" />
                    <RANKING place="22" resultid="928" />
                    <RANKING place="18" resultid="937" />
                    <RANKING place="7" resultid="967" />
                    <RANKING place="21" resultid="1883" />
                    <RANKING place="10" resultid="2026" />
                    <RANKING place="15" resultid="2065" />
                    <RANKING place="13" resultid="3841" />
                    <RANKING place="16" resultid="4187" />
                    <RANKING place="1" resultid="4379" />
                    <RANKING place="3" resultid="4399" />
                    <RANKING place="4" resultid="4496" />
                    <RANKING place="11" resultid="4521" />
                    <RANKING place="6" resultid="4525" />
                    <RANKING place="14" resultid="4682" />
                    <RANKING place="12" resultid="4715" />
                    <RANKING place="8" resultid="4925" />
                    <RANKING place="5" resultid="5018" />
                    <RANKING place="2" resultid="5657" />
                    <RANKING place="20" resultid="6073" />
                    <RANKING place="17" resultid="6106" />
                    <RANKING place="9" resultid="6165" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9" agemax="9" agemin="9" name="Jahrgang 2014">
                  <RANKINGS>
                    <RANKING place="3" resultid="881" />
                    <RANKING place="27" resultid="924" />
                    <RANKING place="34" resultid="979" />
                    <RANKING place="36" resultid="984" />
                    <RANKING place="33" resultid="1007" />
                    <RANKING place="4" resultid="1017" />
                    <RANKING place="8" resultid="1602" />
                    <RANKING place="18" resultid="1619" />
                    <RANKING place="15" resultid="1968" />
                    <RANKING place="17" resultid="2000" />
                    <RANKING place="35" resultid="2018" />
                    <RANKING place="32" resultid="2049" />
                    <RANKING place="2" resultid="2055" />
                    <RANKING place="12" resultid="4035" />
                    <RANKING place="11" resultid="4048" />
                    <RANKING place="20" resultid="4119" />
                    <RANKING place="6" resultid="4144" />
                    <RANKING place="5" resultid="4194" />
                    <RANKING place="10" resultid="4200" />
                    <RANKING place="24" resultid="4208" />
                    <RANKING place="26" resultid="4212" />
                    <RANKING place="7" resultid="4232" />
                    <RANKING place="19" resultid="4239" />
                    <RANKING place="29" resultid="4535" />
                    <RANKING place="14" resultid="4657" />
                    <RANKING place="9" resultid="4772" />
                    <RANKING place="16" resultid="5051" />
                    <RANKING place="25" resultid="5186" />
                    <RANKING place="30" resultid="5198" />
                    <RANKING place="28" resultid="5410" />
                    <RANKING place="31" resultid="5470" />
                    <RANKING place="22" resultid="5602" />
                    <RANKING place="23" resultid="5960" />
                    <RANKING place="13" resultid="6219" />
                    <RANKING place="1" resultid="6244" />
                    <RANKING place="21" resultid="6257" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
          </EVENTS>
        </SESSION>
        <SESSION number="4" date="2023-07-02">
          <EVENTS>
            <EVENT eventid="31" number="31" gender="F" round="TIM">
              <SWIMSTYLE stroke="FLY" name="50 Delphinbeinbewegung Frauen" technique="KICK" relaycount="1" distance="50" />
              <HEATS>
                <HEAT heatid="31001" number="1" />
                <HEAT heatid="31002" number="2" />
                <HEAT heatid="31003" number="3" />
                <HEAT heatid="31004" number="4" />
                <HEAT heatid="31005" number="5" />
                <HEAT heatid="31006" number="6" />
                <HEAT heatid="31007" number="7" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="9" agemax="9" agemin="9" name="Jahrgang 2014">
                  <RANKINGS>
                    <RANKING place="25" resultid="835" />
                    <RANKING place="11" resultid="908" />
                    <RANKING place="9" resultid="919" />
                    <RANKING place="18" resultid="932" />
                    <RANKING place="1" resultid="963" />
                    <RANKING place="8" resultid="1634" />
                    <RANKING place="2" resultid="1639" />
                    <RANKING place="22" resultid="4086" />
                    <RANKING place="6" resultid="4123" />
                    <RANKING place="10" resultid="4277" />
                    <RANKING place="14" resultid="4308" />
                    <RANKING place="3" resultid="4330" />
                    <RANKING place="7" resultid="4335" />
                    <RANKING place="13" resultid="4365" />
                    <RANKING place="15" resultid="4463" />
                    <RANKING place="5" resultid="4768" />
                    <RANKING place="24" resultid="5047" />
                    <RANKING place="16" resultid="5080" />
                    <RANKING place="21" resultid="5104" />
                    <RANKING place="19" resultid="5216" />
                    <RANKING place="12" resultid="5485" />
                    <RANKING place="17" resultid="5555" />
                    <RANKING place="23" resultid="5562" />
                    <RANKING place="20" resultid="5598" />
                    <RANKING place="4" resultid="5680" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1" agemax="10" agemin="10" name="Jahrgang 2013">
                  <RANKINGS>
                    <RANKING place="5" resultid="475" />
                    <RANKING place="10" resultid="779" />
                    <RANKING place="4" resultid="885" />
                    <RANKING place="11" resultid="947" />
                    <RANKING place="13" resultid="3824" />
                    <RANKING place="8" resultid="4359" />
                    <RANKING place="6" resultid="4430" />
                    <RANKING place="1" resultid="4446" />
                    <RANKING place="3" resultid="4512" />
                    <RANKING place="7" resultid="4620" />
                    <RANKING place="12" resultid="4751" />
                    <RANKING place="9" resultid="5099" />
                    <RANKING place="2" resultid="5444" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2" agemax="11" agemin="11" name="Jahrgang 2012">
                  <RANKINGS>
                    <RANKING place="8" resultid="1644" />
                    <RANKING place="3" resultid="4324" />
                    <RANKING place="4" resultid="4915" />
                    <RANKING place="6" resultid="5110" />
                    <RANKING place="5" resultid="5234" />
                    <RANKING place="1" resultid="5345" />
                    <RANKING place="2" resultid="5846" />
                    <RANKING place="7" resultid="6181" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="32" number="32" gender="M" round="TIM">
              <SWIMSTYLE stroke="FLY" name="50 Delphinbeinbewegung Frauen" technique="KICK" relaycount="1" distance="50" />
              <HEATS>
                <HEAT heatid="32001" number="1" />
                <HEAT heatid="32002" number="2" />
                <HEAT heatid="32003" number="3" />
                <HEAT heatid="32004" number="4" />
                <HEAT heatid="32005" number="5" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="9" agemax="9" agemin="9" name="Jahrgang 2014">
                  <RANKINGS>
                    <RANKING place="2" resultid="880" />
                    <RANKING place="8" resultid="1999" />
                    <RANKING place="9" resultid="4036" />
                    <RANKING place="4" resultid="4145" />
                    <RANKING place="3" resultid="4195" />
                    <RANKING place="5" resultid="4233" />
                    <RANKING place="12" resultid="4658" />
                    <RANKING place="6" resultid="4773" />
                    <RANKING place="13" resultid="5052" />
                    <RANKING place="10" resultid="5199" />
                    <RANKING place="11" resultid="5471" />
                    <RANKING place="7" resultid="5603" />
                    <RANKING place="1" resultid="5732" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1" agemax="10" agemin="10" name="Jahrgang 2013">
                  <RANKINGS>
                    <RANKING place="7" resultid="848" />
                    <RANKING place="4" resultid="2129" />
                    <RANKING place="11" resultid="3801" />
                    <RANKING place="9" resultid="3837" />
                    <RANKING place="10" resultid="4043" />
                    <RANKING place="3" resultid="4346" />
                    <RANKING place="1" resultid="4368" />
                    <RANKING place="2" resultid="4423" />
                    <RANKING place="6" resultid="5175" />
                    <RANKING place="8" resultid="5947" />
                    <RANKING place="5" resultid="6264" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2" agemax="11" agemin="11" name="Jahrgang 2012">
                  <RANKINGS>
                    <RANKING place="1" resultid="191" />
                    <RANKING place="6" resultid="997" />
                    <RANKING place="4" resultid="2133" />
                    <RANKING place="3" resultid="4244" />
                    <RANKING place="2" resultid="4402" />
                    <RANKING place="7" resultid="4483" />
                    <RANKING place="5" resultid="6012" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="33" number="33" gender="F" round="TIM">
              <SWIMSTYLE stroke="FREE" relaycount="1" distance="100" />
              <HEATS>
                <HEAT heatid="33001" number="1" />
                <HEAT heatid="33002" number="2" />
                <HEAT heatid="33003" number="3" />
                <HEAT heatid="33004" number="4" />
                <HEAT heatid="33005" number="5" />
                <HEAT heatid="33006" number="6" />
                <HEAT heatid="33007" number="7" />
                <HEAT heatid="33008" number="8" />
                <HEAT heatid="33009" number="9" />
                <HEAT heatid="33010" number="10" />
                <HEAT heatid="33011" number="11" />
                <HEAT heatid="33012" number="12" />
                <HEAT heatid="33013" number="13" />
                <HEAT heatid="33014" number="14" />
                <HEAT heatid="33015" number="15" />
                <HEAT heatid="33016" number="16" />
                <HEAT heatid="33017" number="17" />
                <HEAT heatid="33018" number="18" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="9" agemax="9" agemin="9" name="Jahrgang 2014">
                  <RANKINGS>
                    <RANKING place="5" resultid="800" />
                    <RANKING place="14" resultid="907" />
                    <RANKING place="2" resultid="962" />
                    <RANKING place="7" resultid="1655" />
                    <RANKING place="10" resultid="1659" />
                    <RANKING place="9" resultid="1905" />
                    <RANKING place="18" resultid="2013" />
                    <RANKING place="19" resultid="2093" />
                    <RANKING place="12" resultid="4087" />
                    <RANKING place="21" resultid="4096" />
                    <RANKING place="11" resultid="4124" />
                    <RANKING place="1" resultid="4282" />
                    <RANKING place="17" resultid="4313" />
                    <RANKING place="4" resultid="4383" />
                    <RANKING place="8" resultid="4412" />
                    <RANKING place="3" resultid="4435" />
                    <RANKING place="20" resultid="5023" />
                    <RANKING place="16" resultid="5028" />
                    <RANKING place="13" resultid="5048" />
                    <RANKING place="6" resultid="5081" />
                    <RANKING place="15" resultid="5116" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1" agemax="10" agemin="10" name="Jahrgang 2013">
                  <RANKINGS>
                    <RANKING place="6" resultid="12" />
                    <RANKING place="7" resultid="476" />
                    <RANKING place="11" resultid="761" />
                    <RANKING place="17" resultid="778" />
                    <RANKING place="12" resultid="1917" />
                    <RANKING place="20" resultid="1963" />
                    <RANKING place="19" resultid="1995" />
                    <RANKING place="18" resultid="3727" />
                    <RANKING place="16" resultid="4356" />
                    <RANKING place="14" resultid="4360" />
                    <RANKING place="4" resultid="4475" />
                    <RANKING place="2" resultid="4516" />
                    <RANKING place="13" resultid="4752" />
                    <RANKING place="1" resultid="5144" />
                    <RANKING place="8" resultid="5194" />
                    <RANKING place="15" resultid="5250" />
                    <RANKING place="10" resultid="5479" />
                    <RANKING place="3" resultid="5578" />
                    <RANKING place="9" resultid="5833" />
                    <RANKING place="5" resultid="6109" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2" agemax="11" agemin="11" name="Jahrgang 2012">
                  <RANKINGS>
                    <RANKING place="4" resultid="20" />
                    <RANKING place="6" resultid="183" />
                    <RANKING place="9" resultid="805" />
                    <RANKING place="1" resultid="955" />
                    <RANKING place="7" resultid="1612" />
                    <RANKING place="17" resultid="1649" />
                    <RANKING place="16" resultid="3810" />
                    <RANKING place="8" resultid="4325" />
                    <RANKING place="12" resultid="4862" />
                    <RANKING place="23" resultid="4876" />
                    <RANKING place="19" resultid="5039" />
                    <RANKING place="15" resultid="5111" />
                    <RANKING place="5" resultid="5182" />
                    <RANKING place="18" resultid="5495" />
                    <RANKING place="22" resultid="5614" />
                    <RANKING place="24" resultid="5622" />
                    <RANKING place="3" resultid="5640" />
                    <RANKING place="13" resultid="5647" />
                    <RANKING place="20" resultid="5675" />
                    <RANKING place="2" resultid="5715" />
                    <RANKING place="14" resultid="5724" />
                    <RANKING place="25" resultid="5820" />
                    <RANKING place="21" resultid="5976" />
                    <RANKING place="11" resultid="6039" />
                    <RANKING place="10" resultid="6236" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="13" agemin="12" name="Jahrgang 2010/2011">
                  <RANKINGS>
                    <RANKING place="13" resultid="23" />
                    <RANKING place="5" resultid="135" />
                    <RANKING place="28" resultid="151" />
                    <RANKING place="9" resultid="159" />
                    <RANKING place="3" resultid="175" />
                    <RANKING place="2" resultid="615" />
                    <RANKING place="8" resultid="972" />
                    <RANKING place="17" resultid="1914" />
                    <RANKING place="14" resultid="1944" />
                    <RANKING place="22" resultid="2032" />
                    <RANKING place="34" resultid="2098" />
                    <RANKING place="29" resultid="2102" />
                    <RANKING place="4" resultid="2137" />
                    <RANKING place="35" resultid="3739" />
                    <RANKING place="36" resultid="3752" />
                    <RANKING place="23" resultid="3772" />
                    <RANKING place="11" resultid="3845" />
                    <RANKING place="32" resultid="4303" />
                    <RANKING place="30" resultid="4699" />
                    <RANKING place="24" resultid="4848" />
                    <RANKING place="15" resultid="4869" />
                    <RANKING place="25" resultid="4883" />
                    <RANKING place="18" resultid="4932" />
                    <RANKING place="16" resultid="4935" />
                    <RANKING place="33" resultid="5004" />
                    <RANKING place="21" resultid="5032" />
                    <RANKING place="27" resultid="5088" />
                    <RANKING place="26" resultid="5150" />
                    <RANKING place="12" resultid="5152" />
                    <RANKING place="19" resultid="5211" />
                    <RANKING place="7" resultid="5242" />
                    <RANKING place="9" resultid="5299" />
                    <RANKING place="1" resultid="5502" />
                    <RANKING place="31" resultid="5764" />
                    <RANKING place="20" resultid="5792" />
                    <RANKING place="6" resultid="6115" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6" agemax="15" agemin="14" name="Jahrgang 2008/2009">
                  <RANKINGS>
                    <RANKING place="1" resultid="610" />
                    <RANKING place="20" resultid="1922" />
                    <RANKING place="14" resultid="4292" />
                    <RANKING place="3" resultid="4584" />
                    <RANKING place="7" resultid="4889" />
                    <RANKING place="11" resultid="4945" />
                    <RANKING place="17" resultid="4965" />
                    <RANKING place="4" resultid="4997" />
                    <RANKING place="8" resultid="5276" />
                    <RANKING place="19" resultid="5296" />
                    <RANKING place="10" resultid="5333" />
                    <RANKING place="2" resultid="5357" />
                    <RANKING place="5" resultid="5434" />
                    <RANKING place="9" resultid="5611" />
                    <RANKING place="16" resultid="5737" />
                    <RANKING place="15" resultid="5876" />
                    <RANKING place="12" resultid="5916" />
                    <RANKING place="13" resultid="5964" />
                    <RANKING place="18" resultid="6191" />
                    <RANKING place="6" resultid="6363" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8" agemax="17" agemin="16" name="Jahrgang 2006/2007">
                  <RANKINGS>
                    <RANKING place="5" resultid="3725" />
                    <RANKING place="8" resultid="3744" />
                    <RANKING place="6" resultid="4653" />
                    <RANKING place="3" resultid="4704" />
                    <RANKING place="4" resultid="4842" />
                    <RANKING place="7" resultid="4962" />
                    <RANKING place="2" resultid="4968" />
                    <RANKING place="9" resultid="4977" />
                    <RANKING place="1" resultid="5489" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="34" number="34" gender="M" round="TIM">
              <SWIMSTYLE stroke="FREE" relaycount="1" distance="100" />
              <HEATS>
                <HEAT heatid="34001" number="1" />
                <HEAT heatid="34002" number="2" />
                <HEAT heatid="34003" number="3" />
                <HEAT heatid="34004" number="4" />
                <HEAT heatid="34005" number="5" />
                <HEAT heatid="34006" number="6" />
                <HEAT heatid="34007" number="7" />
                <HEAT heatid="34008" number="8" />
                <HEAT heatid="34009" number="9" />
                <HEAT heatid="34010" number="10" />
                <HEAT heatid="34011" number="11" />
                <HEAT heatid="34012" number="12" />
                <HEAT heatid="34013" number="13" />
                <HEAT heatid="34014" number="14" />
                <HEAT heatid="34015" number="15" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="9" agemax="9" agemin="9" name="Jahrgang 2014">
                  <RANKINGS>
                    <RANKING place="2" resultid="1016" />
                    <RANKING place="5" resultid="1601" />
                    <RANKING place="7" resultid="1618" />
                    <RANKING place="6" resultid="1967" />
                    <RANKING place="1" resultid="2054" />
                    <RANKING place="3" resultid="4049" />
                    <RANKING place="9" resultid="4146" />
                    <RANKING place="4" resultid="5053" />
                    <RANKING place="8" resultid="5187" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1" agemax="10" agemin="10" name="Jahrgang 2013">
                  <RANKINGS>
                    <RANKING place="16" resultid="758" />
                    <RANKING place="12" resultid="847" />
                    <RANKING place="4" resultid="942" />
                    <RANKING place="22" resultid="2034" />
                    <RANKING place="1" resultid="3434" />
                    <RANKING place="24" resultid="3735" />
                    <RANKING place="25" resultid="3800" />
                    <RANKING place="7" resultid="4044" />
                    <RANKING place="6" resultid="4054" />
                    <RANKING place="19" resultid="4102" />
                    <RANKING place="10" resultid="4179" />
                    <RANKING place="14" resultid="4369" />
                    <RANKING place="3" resultid="4394" />
                    <RANKING place="11" resultid="4764" />
                    <RANKING place="21" resultid="4780" />
                    <RANKING place="8" resultid="4987" />
                    <RANKING place="23" resultid="5067" />
                    <RANKING place="20" resultid="5176" />
                    <RANKING place="15" resultid="5540" />
                    <RANKING place="18" resultid="5591" />
                    <RANKING place="5" resultid="5628" />
                    <RANKING place="9" resultid="5839" />
                    <RANKING place="17" resultid="5892" />
                    <RANKING place="2" resultid="5955" />
                    <RANKING place="13" resultid="6202" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2" agemax="11" agemin="11" name="Jahrgang 2012">
                  <RANKINGS>
                    <RANKING place="2" resultid="127" />
                    <RANKING place="27" resultid="168" />
                    <RANKING place="1" resultid="192" />
                    <RANKING place="18" resultid="782" />
                    <RANKING place="5" resultid="818" />
                    <RANKING place="21" resultid="855" />
                    <RANKING place="9" resultid="913" />
                    <RANKING place="20" resultid="989" />
                    <RANKING place="23" resultid="996" />
                    <RANKING place="8" resultid="2005" />
                    <RANKING place="7" resultid="3455" />
                    <RANKING place="28" resultid="3746" />
                    <RANKING place="13" resultid="4070" />
                    <RANKING place="12" resultid="4245" />
                    <RANKING place="10" resultid="4272" />
                    <RANKING place="15" resultid="4419" />
                    <RANKING place="6" resultid="4453" />
                    <RANKING place="26" resultid="4484" />
                    <RANKING place="16" resultid="4721" />
                    <RANKING place="14" resultid="4800" />
                    <RANKING place="19" resultid="4830" />
                    <RANKING place="3" resultid="5522" />
                    <RANKING place="17" resultid="5529" />
                    <RANKING place="22" resultid="5571" />
                    <RANKING place="4" resultid="5691" />
                    <RANKING place="25" resultid="5854" />
                    <RANKING place="11" resultid="5943" />
                    <RANKING place="24" resultid="6013" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="13" agemin="12" name="Jahrgang 2010/2011">
                  <RANKINGS>
                    <RANKING place="6" resultid="119" />
                    <RANKING place="7" resultid="143" />
                    <RANKING place="3" resultid="768" />
                    <RANKING place="5" resultid="790" />
                    <RANKING place="1" resultid="808" />
                    <RANKING place="20" resultid="1887" />
                    <RANKING place="13" resultid="1936" />
                    <RANKING place="14" resultid="1983" />
                    <RANKING place="19" resultid="2045" />
                    <RANKING place="15" resultid="2088" />
                    <RANKING place="9" resultid="3440" />
                    <RANKING place="18" resultid="3732" />
                    <RANKING place="11" resultid="4289" />
                    <RANKING place="4" resultid="4631" />
                    <RANKING place="10" resultid="4896" />
                    <RANKING place="12" resultid="4991" />
                    <RANKING place="8" resultid="5246" />
                    <RANKING place="17" resultid="5268" />
                    <RANKING place="2" resultid="5700" />
                    <RANKING place="16" resultid="6168" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6" agemax="15" agemin="14" name="Jahrgang 2008/2009">
                  <RANKINGS>
                    <RANKING place="14" resultid="3713" />
                    <RANKING place="17" resultid="3768" />
                    <RANKING place="12" resultid="4265" />
                    <RANKING place="4" resultid="4319" />
                    <RANKING place="6" resultid="4664" />
                    <RANKING place="7" resultid="4785" />
                    <RANKING place="13" resultid="4809" />
                    <RANKING place="15" resultid="4823" />
                    <RANKING place="5" resultid="4855" />
                    <RANKING place="9" resultid="4909" />
                    <RANKING place="8" resultid="4954" />
                    <RANKING place="10" resultid="5071" />
                    <RANKING place="16" resultid="5430" />
                    <RANKING place="1" resultid="5511" />
                    <RANKING place="2" resultid="5903" />
                    <RANKING place="3" resultid="6001" />
                    <RANKING place="11" resultid="6098" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8" agemax="17" agemin="16" name="Jahrgang 2006/2007">
                  <RANKINGS>
                    <RANKING place="4" resultid="3482" />
                    <RANKING place="8" resultid="3796" />
                    <RANKING place="1" resultid="4710" />
                    <RANKING place="6" resultid="4836" />
                    <RANKING place="3" resultid="5137" />
                    <RANKING place="2" resultid="5317" />
                    <RANKING place="7" resultid="5374" />
                    <RANKING place="5" resultid="5583" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="35" number="35" gender="F" round="TIM">
              <SWIMSTYLE stroke="FLY" relaycount="1" distance="100" />
              <HEATS>
                <HEAT heatid="35001" number="1" />
                <HEAT heatid="35002" number="2" />
                <HEAT heatid="35003" number="3" />
                <HEAT heatid="35004" number="4" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="10" agemin="10" name="Jahrgang 2013">
                  <RANKINGS>
                    <RANKING place="1" resultid="764" />
                    <RANKING place="2" resultid="797" />
                    <RANKING place="3" resultid="4447" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2" agemax="11" agemin="11" name="Jahrgang 2012">
                  <RANKINGS>
                    <RANKING place="2" resultid="1954" />
                    <RANKING place="4" resultid="4480" />
                    <RANKING place="5" resultid="4922" />
                    <RANKING place="3" resultid="5235" />
                    <RANKING place="1" resultid="5346" />
                    <RANKING place="6" resultid="5935" />
                    <RANKING place="7" resultid="6028" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="13" agemin="12" name="Jahrgang 2010/2011">
                  <RANKINGS>
                    <RANKING place="2" resultid="136" />
                    <RANKING place="5" resultid="152" />
                    <RANKING place="1" resultid="176" />
                    <RANKING place="4" resultid="5153" />
                    <RANKING place="3" resultid="5406" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6" agemax="15" agemin="14" name="Jahrgang 2008/2009">
                  <RANKINGS>
                    <RANKING place="7" resultid="3720" />
                    <RANKING place="4" resultid="3820" />
                    <RANKING place="5" resultid="4998" />
                    <RANKING place="2" resultid="5358" />
                    <RANKING place="6" resultid="5667" />
                    <RANKING place="1" resultid="5878" />
                    <RANKING place="3" resultid="6277" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8" agemax="17" agemin="16" name="Jahrgang 2006/2007">
                  <RANKINGS>
                    <RANKING place="3" resultid="3808" />
                    <RANKING place="2" resultid="4705" />
                    <RANKING place="1" resultid="4732" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="36" number="36" gender="M" round="TIM">
              <SWIMSTYLE stroke="FLY" relaycount="1" distance="100" />
              <HEATS>
                <HEAT heatid="36001" number="1" />
                <HEAT heatid="36002" number="2" />
                <HEAT heatid="36003" number="3" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="10" agemin="10" name="Jahrgang 2013">
                  <RANKINGS>
                    <RANKING place="4" resultid="2128" />
                    <RANKING place="1" resultid="4347" />
                    <RANKING place="2" resultid="5629" />
                    <RANKING place="3" resultid="5840" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2" agemax="11" agemin="11" name="Jahrgang 2012">
                  <RANKINGS>
                    <RANKING place="3" resultid="2132" />
                    <RANKING place="2" resultid="4403" />
                    <RANKING place="4" resultid="5311" />
                    <RANKING place="1" resultid="6186" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="13" agemin="12" name="Jahrgang 2010/2011">
                  <RANKINGS>
                    <RANKING place="3" resultid="767" />
                    <RANKING place="2" resultid="789" />
                    <RANKING place="1" resultid="869" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6" agemax="15" agemin="14" name="Jahrgang 2008/2009">
                  <RANKINGS>
                    <RANKING place="4" resultid="3816" />
                    <RANKING place="3" resultid="4955" />
                    <RANKING place="2" resultid="5364" />
                    <RANKING place="1" resultid="6020" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8" agemax="17" agemin="16" name="Jahrgang 2006/2007">
                  <RANKINGS>
                    <RANKING place="1" resultid="5138" />
                    <RANKING place="2" resultid="5375" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="37" number="37" gender="F" round="TIM">
              <SWIMSTYLE stroke="BACK" relaycount="1" distance="200" />
              <HEATS>
                <HEAT heatid="37001" number="1" />
                <HEAT heatid="37002" number="2" />
                <HEAT heatid="37003" number="3" />
                <HEAT heatid="37004" number="4" />
                <HEAT heatid="37005" number="5" />
                <HEAT heatid="37006" number="6" />
                <HEAT heatid="37007" number="7" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="10" agemin="10" name="Jahrgang 2013">
                  <RANKINGS>
                    <RANKING place="4" resultid="13" />
                    <RANKING place="7" resultid="1916" />
                    <RANKING place="3" resultid="4458" />
                    <RANKING place="6" resultid="4476" />
                    <RANKING place="2" resultid="4513" />
                    <RANKING place="8" resultid="4517" />
                    <RANKING place="1" resultid="5445" />
                    <RANKING place="9" resultid="5480" />
                    <RANKING place="10" resultid="6053" />
                    <RANKING place="5" resultid="6110" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2" agemax="11" agemin="11" name="Jahrgang 2012">
                  <RANKINGS>
                    <RANKING place="8" resultid="184" />
                    <RANKING place="9" resultid="804" />
                    <RANKING place="11" resultid="954" />
                    <RANKING place="12" resultid="1595" />
                    <RANKING place="5" resultid="1990" />
                    <RANKING place="3" resultid="4509" />
                    <RANKING place="6" resultid="4916" />
                    <RANKING place="10" resultid="5648" />
                    <RANKING place="1" resultid="5716" />
                    <RANKING place="2" resultid="5847" />
                    <RANKING place="13" resultid="5936" />
                    <RANKING place="7" resultid="6040" />
                    <RANKING place="14" resultid="6182" />
                    <RANKING place="4" resultid="6237" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="13" agemin="12" name="Jahrgang 2010/2011">
                  <RANKINGS>
                    <RANKING place="10" resultid="24" />
                    <RANKING place="5" resultid="160" />
                    <RANKING place="6" resultid="219" />
                    <RANKING place="3" resultid="971" />
                    <RANKING place="13" resultid="1913" />
                    <RANKING place="11" resultid="1985" />
                    <RANKING place="12" resultid="2031" />
                    <RANKING place="9" resultid="2059" />
                    <RANKING place="4" resultid="2136" />
                    <RANKING place="8" resultid="4936" />
                    <RANKING place="7" resultid="5300" />
                    <RANKING place="2" resultid="5395" />
                    <RANKING place="14" resultid="5765" />
                    <RANKING place="1" resultid="6116" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6" agemax="15" agemin="14" name="Jahrgang 2008/2009">
                  <RANKINGS>
                    <RANKING place="1" resultid="2010" />
                    <RANKING place="3" resultid="5277" />
                    <RANKING place="2" resultid="5334" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8" agemax="17" agemin="16" name="Jahrgang 2006/2007" />
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="38" number="38" gender="M" round="TIM">
              <SWIMSTYLE stroke="BACK" relaycount="1" distance="200" />
              <HEATS>
                <HEAT heatid="38001" number="1" />
                <HEAT heatid="38002" number="2" />
                <HEAT heatid="38003" number="3" />
                <HEAT heatid="38004" number="4" />
                <HEAT heatid="38005" number="5" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="10" agemin="10" name="Jahrgang 2013">
                  <RANKINGS>
                    <RANKING place="1" resultid="941" />
                    <RANKING place="5" resultid="1628" />
                    <RANKING place="9" resultid="4424" />
                    <RANKING place="3" resultid="4500" />
                    <RANKING place="8" resultid="5541" />
                    <RANKING place="6" resultid="5893" />
                    <RANKING place="2" resultid="5948" />
                    <RANKING place="4" resultid="5956" />
                    <RANKING place="7" resultid="6265" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2" agemax="11" agemin="11" name="Jahrgang 2012">
                  <RANKINGS>
                    <RANKING place="1" resultid="128" />
                    <RANKING place="2" resultid="817" />
                    <RANKING place="10" resultid="854" />
                    <RANKING place="8" resultid="912" />
                    <RANKING place="9" resultid="988" />
                    <RANKING place="5" resultid="2004" />
                    <RANKING place="7" resultid="4420" />
                    <RANKING place="6" resultid="4454" />
                    <RANKING place="11" resultid="5312" />
                    <RANKING place="4" resultid="5530" />
                    <RANKING place="3" resultid="5944" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="13" agemin="12" name="Jahrgang 2010/2011">
                  <RANKINGS>
                    <RANKING place="2" resultid="120" />
                    <RANKING place="3" resultid="144" />
                    <RANKING place="1" resultid="807" />
                    <RANKING place="6" resultid="1929" />
                    <RANKING place="5" resultid="1935" />
                    <RANKING place="8" resultid="1982" />
                    <RANKING place="7" resultid="2087" />
                    <RANKING place="9" resultid="5269" />
                    <RANKING place="4" resultid="5752" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6" agemax="15" agemin="14" name="Jahrgang 2008/2009">
                  <RANKINGS>
                    <RANKING place="2" resultid="4786" />
                    <RANKING place="1" resultid="5388" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8" agemax="17" agemin="16" name="Jahrgang 2006/2007">
                  <RANKINGS>
                    <RANKING place="2" resultid="3783" />
                    <RANKING place="3" resultid="4711" />
                    <RANKING place="1" resultid="5318" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
          </EVENTS>
        </SESSION>
      </SESSIONS>
      <CLUBS>
        <CLUB name="1. Chemnitzer Tauchverein e.V." nation="GER" region="20" code="0">
          <ATHLETES>
            <ATHLETE athleteid="447" birthdate="2012-01-01" gender="M" lastname="Ilianyi" firstname="Yan" license="0">
              <RESULTS>
                <RESULT resultid="2156" eventid="40" swimtime="00:02:54.16" lane="5" heatid="40001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:22.17" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="2155" eventid="46" swimtime="00:01:22.77" lane="3" heatid="46001" />
                <RESULT resultid="2154" eventid="50" swimtime="00:00:32.47" lane="3" heatid="50002" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="448" birthdate="2010-01-01" gender="M" lastname="Yemelianov" firstname="Viktor" license="0">
              <RESULTS>
                <RESULT resultid="2159" eventid="40" swimtime="00:02:30.71" lane="6" heatid="40001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:10.23" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="2158" eventid="46" swimtime="00:01:07.38" lane="8" heatid="46001" />
                <RESULT resultid="2157" eventid="50" swimtime="00:00:28.90" lane="6" heatid="50001" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="449" birthdate="2010-01-01" gender="F" lastname="Bluhm" firstname="Suna" license="0">
              <RESULTS>
                <RESULT resultid="2162" eventid="41" swimtime="00:00:13.62" lane="3" heatid="41002" />
                <RESULT resultid="2161" eventid="45" swimtime="00:01:03.73" lane="1" heatid="45005" />
                <RESULT resultid="2160" eventid="49" swimtime="00:00:28.61" lane="1" heatid="49004" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="450" birthdate="2009-01-01" gender="M" lastname="Elle" firstname="Simon" license="0">
              <RESULTS>
                <RESULT resultid="2166" eventid="42" swimtime="00:00:16.87" lane="7" heatid="42002" />
                <RESULT resultid="2165" eventid="46" swimtime="00:01:13.70" lane="2" heatid="46002" />
                <RESULT resultid="2164" eventid="48" swimtime="00:00:40.33" lane="6" heatid="48001" />
                <RESULT resultid="2163" eventid="50" swimtime="00:00:33.28" lane="5" heatid="50002" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="451" birthdate="2012-01-01" gender="F" lastname="Gralka" firstname="Lilou" license="0">
              <RESULTS>
                <RESULT resultid="2168" eventid="45" swimtime="00:01:23.02" lane="3" heatid="45001" />
                <RESULT resultid="2167" eventid="49" swimtime="00:00:35.93" lane="2" heatid="49001" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="452" birthdate="2007-01-01" gender="F" lastname="Ullrich" firstname="Johanna Hermine" license="0">
              <RESULTS>
                <RESULT resultid="2172" eventid="39" status="DNS" swimtime="00:00:00.00" lane="5" heatid="39003" />
                <RESULT resultid="2171" eventid="41" swimtime="00:00:13.14" lane="8" heatid="41005" />
                <RESULT resultid="2170" eventid="45" swimtime="00:00:56.14" lane="6" heatid="45006" />
                <RESULT resultid="2169" eventid="49" swimtime="00:00:25.01" lane="7" heatid="49005" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="453" birthdate="2008-01-01" gender="F" lastname="Franke" firstname="Jenny" license="0">
              <RESULTS>
                <RESULT resultid="2176" eventid="39" swimtime="00:01:53.22" lane="3" heatid="39003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:54.09" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="2175" eventid="41" swimtime="00:00:10.96" lane="7" heatid="41005" />
                <RESULT resultid="2174" eventid="45" swimtime="00:00:48.08" lane="5" heatid="45006" />
                <RESULT resultid="2173" eventid="49" swimtime="00:00:21.74" lane="2" heatid="49005" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="454" birthdate="2012-01-01" gender="F" lastname="Laasner" firstname="Ida Marie" license="0">
              <RESULTS>
                <RESULT resultid="2178" eventid="45" swimtime="00:01:25.43" lane="5" heatid="45001" />
                <RESULT resultid="2177" eventid="49" swimtime="00:00:35.78" lane="7" heatid="49001" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="455" birthdate="2010-01-01" gender="F" lastname="Siegert" firstname="Emilia" license="0">
              <RESULTS>
                <RESULT resultid="2182" eventid="39" swimtime="00:02:15.99" lane="4" heatid="39002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:05.06" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="2181" eventid="41" swimtime="00:00:14.10" lane="5" heatid="41002" />
                <RESULT resultid="2180" eventid="45" swimtime="00:00:59.84" lane="7" heatid="45005" />
                <RESULT resultid="2179" eventid="49" swimtime="00:00:26.91" lane="8" heatid="49004" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="456" birthdate="2006-01-01" gender="M" lastname="Lorenz" firstname="Emil" license="0">
              <RESULTS>
                <RESULT resultid="2186" eventid="42" swimtime="00:00:09.18" lane="3" heatid="42003" />
                <RESULT resultid="2185" eventid="46" swimtime="00:00:43.33" lane="3" heatid="46003" />
                <RESULT resultid="2184" eventid="48" swimtime="00:00:24.94" lane="5" heatid="48001" />
                <RESULT resultid="2183" eventid="50" swimtime="00:00:19.18" lane="4" heatid="50003" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="457" birthdate="2013-01-01" gender="M" lastname="Schiller" firstname="Ben" license="0">
              <RESULTS>
                <RESULT resultid="2189" eventid="40" swimtime="00:03:17.97" lane="3" heatid="40001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:32.95" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="2188" eventid="46" swimtime="00:01:34.40" lane="4" heatid="46001" />
                <RESULT resultid="2187" eventid="50" swimtime="00:00:40.65" lane="1" heatid="50002" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="458" birthdate="2009-01-01" gender="M" lastname="Müller" firstname="Alwin" license="0">
              <RESULTS>
                <RESULT resultid="2193" eventid="40" swimtime="00:02:12.76" lane="2" heatid="40002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:02.27" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="2192" eventid="42" swimtime="00:00:15.88" lane="8" heatid="42003" />
                <RESULT resultid="2191" eventid="46" swimtime="00:01:00.26" lane="8" heatid="46003" />
                <RESULT resultid="2190" eventid="50" status="DNS" swimtime="00:00:00.00" lane="4" heatid="50002" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="891" birthdate="2011-01-01" gender="F" lastname="Nisch" firstname="Hanna Maria" license="0">
              <RESULTS>
                <RESULT resultid="4180" eventid="39" swimtime="00:02:13.96" lane="5" heatid="39002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:05.61" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="4181" eventid="41" swimtime="00:00:13.41" lane="1" heatid="41004" />
                <RESULT resultid="4182" eventid="45" swimtime="00:00:58.10" lane="3" heatid="45005" />
                <RESULT resultid="4183" eventid="49" swimtime="00:00:26.14" lane="2" heatid="49004" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="ATSV Freiberg e.V." nation="GER" region="12" code="3324">
          <ATHLETES>
            <ATHLETE athleteid="905" birthdate="2014-01-01" gender="M" lastname="Kiekebelt" firstname="Alexander" license="445951">
              <RESULTS>
                <RESULT resultid="4235" eventid="18" swimtime="00:01:04.93" lane="2" heatid="18007" />
                <RESULT resultid="4236" eventid="20" swimtime="00:01:01.75" lane="5" heatid="20003" />
                <RESULT resultid="4237" eventid="22" swimtime="00:01:02.02" lane="6" heatid="22005" />
                <RESULT resultid="4238" eventid="26" swimtime="00:00:52.70" lane="3" heatid="26007" />
                <RESULT resultid="4239" eventid="30" swimtime="00:00:46.12" lane="1" heatid="30007" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="906" birthdate="2012-01-01" gender="M" lastname="Tanneberger" firstname="Arian" license="434981">
              <RESULTS>
                <RESULT resultid="4240" eventid="4" swimtime="00:01:48.74" lane="1" heatid="4005" />
                <RESULT resultid="4241" eventid="6" swimtime="00:00:42.22" lane="4" heatid="6005" />
                <RESULT resultid="4242" eventid="22" swimtime="00:00:45.16" lane="6" heatid="22011" />
                <RESULT resultid="4243" eventid="28" swimtime="00:00:55.74" lane="6" heatid="28005" />
                <RESULT resultid="4244" eventid="32" swimtime="00:00:50.66" lane="5" heatid="32004" />
                <RESULT resultid="4245" eventid="34" swimtime="00:01:19.13" lane="1" heatid="34009" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="907" birthdate="2013-01-01" gender="M" lastname="Oehme" firstname="Arvid" license="445060">
              <RESULTS>
                <RESULT resultid="4246" eventid="6" swimtime="00:00:47.52" lane="2" heatid="6002" />
                <RESULT resultid="4247" eventid="11" swimtime="00:01:50.83" lane="2" heatid="11002" />
                <RESULT resultid="4248" eventid="13" swimtime="00:00:38.33" lane="3" heatid="13004" />
                <RESULT resultid="4249" eventid="20" swimtime="00:00:54.67" lane="8" heatid="20007" />
                <RESULT resultid="4250" eventid="24" swimtime="00:03:15.84" lane="7" heatid="24002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:33.70" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="908" birthdate="2015-01-01" gender="F" lastname="Heinz" firstname="Elizabeth" license="471931">
              <RESULTS>
                <RESULT resultid="4251" eventid="19" swimtime="00:01:05.56" lane="4" heatid="19006" />
                <RESULT resultid="4252" eventid="21" swimtime="00:01:08.09" lane="3" heatid="21004" />
                <RESULT resultid="4253" eventid="25" swimtime="00:00:58.54" lane="3" heatid="25005" />
                <RESULT resultid="4254" eventid="27" swimtime="00:01:11.53" lane="5" heatid="27001" />
                <RESULT resultid="4255" eventid="29" swimtime="00:00:54.76" lane="3" heatid="29004" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="909" birthdate="2013-01-01" gender="F" lastname="Queck" firstname="Fabienne" license="451852">
              <RESULTS>
                <RESULT resultid="4256" eventid="3" swimtime="00:02:05.94" lane="4" heatid="3001" />
                <RESULT resultid="4257" eventid="12" swimtime="00:00:48.94" lane="3" heatid="12001" />
                <RESULT resultid="4258" eventid="14" swimtime="00:04:33.56" lane="8" heatid="14002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:02:13.45" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="910" birthdate="2013-01-01" gender="F" lastname="Brocke" firstname="Fiene" license="445947">
              <RESULTS>
                <RESULT resultid="4259" eventid="3" swimtime="00:02:00.32" lane="3" heatid="3002" />
                <RESULT resultid="4260" eventid="5" swimtime="00:00:55.88" lane="6" heatid="5002" />
                <RESULT resultid="4261" eventid="10" swimtime="00:01:57.88" lane="7" heatid="10003" />
                <RESULT resultid="4262" eventid="12" swimtime="00:00:44.46" lane="7" heatid="12002" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="911" birthdate="2008-01-01" gender="M" lastname="Belger" firstname="Finnian" license="364362">
              <RESULTS>
                <RESULT resultid="4263" eventid="20" swimtime="00:00:40.01" lane="2" heatid="20019" />
                <RESULT resultid="4264" eventid="26" swimtime="00:00:41.04" lane="5" heatid="26018" />
                <RESULT resultid="4265" eventid="34" swimtime="00:01:14.72" lane="1" heatid="34011" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="912" birthdate="2012-01-01" gender="M" lastname="Schubert" firstname="Fritz" license="422021">
              <RESULTS>
                <RESULT resultid="4266" eventid="6" swimtime="00:00:45.83" lane="8" heatid="6003" />
                <RESULT resultid="4267" eventid="11" swimtime="00:01:36.12" lane="5" heatid="11005" />
                <RESULT resultid="4268" eventid="13" swimtime="00:00:34.42" lane="6" heatid="13006" />
                <RESULT resultid="4269" eventid="18" swimtime="00:01:00.58" lane="2" heatid="18009" />
                <RESULT resultid="4270" eventid="22" swimtime="00:00:50.87" lane="7" heatid="22011" />
                <RESULT resultid="4271" eventid="26" swimtime="00:00:43.45" lane="8" heatid="26013" />
                <RESULT resultid="4272" eventid="34" swimtime="00:01:17.58" lane="2" heatid="34008" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="913" birthdate="2014-01-01" gender="F" lastname="Ferkinghoff" firstname="Helene" license="445062">
              <RESULTS>
                <RESULT resultid="4273" eventid="17" swimtime="00:01:01.92" lane="3" heatid="17011" />
                <RESULT resultid="4274" eventid="21" swimtime="00:00:55.83" lane="3" heatid="21011" />
                <RESULT resultid="4275" eventid="25" swimtime="00:00:54.73" lane="7" heatid="25011" />
                <RESULT resultid="4276" eventid="29" swimtime="00:00:42.42" lane="2" heatid="29008" />
                <RESULT resultid="4277" eventid="31" swimtime="00:01:03.15" lane="5" heatid="31004" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="914" birthdate="2014-01-01" gender="F" lastname="Riedel" firstname="Hely Margo" license="445061">
              <RESULTS>
                <RESULT resultid="4278" eventid="19" swimtime="00:00:43.86" lane="1" heatid="19021" />
                <RESULT resultid="4279" eventid="25" swimtime="00:00:41.03" lane="8" heatid="25022" />
                <RESULT resultid="4280" eventid="27" swimtime="00:00:54.19" lane="4" heatid="27012" />
                <RESULT resultid="4281" eventid="29" swimtime="00:00:35.44" lane="6" heatid="29013" />
                <RESULT resultid="4282" eventid="33" swimtime="00:01:19.65" lane="2" heatid="33012" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="915" birthdate="2010-01-01" gender="M" lastname="Tanneberger" firstname="Janis" license="407515">
              <RESULTS>
                <RESULT resultid="4283" eventid="4" swimtime="00:01:34.91" lane="8" heatid="4007" />
                <RESULT resultid="4284" eventid="6" swimtime="00:00:38.03" lane="2" heatid="6006" />
                <RESULT resultid="4285" eventid="13" swimtime="00:00:32.71" lane="3" heatid="13011" />
                <RESULT resultid="4286" eventid="15" status="DSQ" swimtime="00:03:32.59" lane="7" heatid="15005" comment="Anschlag bei der 2. Wende erfolgte nicht mir beiden Händen gleichzeitig.">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:43.22" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="4287" eventid="20" swimtime="00:00:43.19" lane="1" heatid="20015" />
                <RESULT resultid="4288" eventid="26" swimtime="00:00:39.66" lane="4" heatid="26019" />
                <RESULT resultid="4289" eventid="34" swimtime="00:01:16.04" lane="5" heatid="34009" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="916" birthdate="2009-01-01" gender="F" lastname="Schierz" firstname="Johanna" license="383730">
              <RESULTS>
                <RESULT resultid="4290" eventid="19" swimtime="00:00:45.41" lane="5" heatid="19023" />
                <RESULT resultid="4291" eventid="25" swimtime="00:00:36.03" lane="2" heatid="25025" />
                <RESULT resultid="4292" eventid="33" swimtime="00:01:12.94" lane="2" heatid="33013" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="917" birthdate="2007-01-01" gender="M" lastname="Frisch" firstname="Jonathan" license="384470">
              <RESULTS>
                <RESULT resultid="4293" eventid="4" swimtime="00:01:24.67" lane="8" heatid="4009" />
                <RESULT resultid="4294" eventid="6" swimtime="00:00:38.49" lane="2" heatid="6005" />
                <RESULT resultid="4295" eventid="13" swimtime="00:00:30.58" lane="1" heatid="13014" />
                <RESULT resultid="4296" eventid="15" swimtime="00:03:09.20" lane="7" heatid="15006">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:30.00" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="4297" eventid="20" swimtime="00:00:38.06" lane="3" heatid="20020" />
                <RESULT resultid="4298" eventid="24" swimtime="00:02:41.38" lane="5" heatid="24006">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:14.99" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="918" birthdate="2013-01-01" gender="F" lastname="Müller" firstname="Lara" license="431998">
              <RESULTS>
                <RESULT resultid="4299" eventid="17" swimtime="00:01:16.20" lane="6" heatid="17008" />
                <RESULT resultid="4300" eventid="21" swimtime="00:01:08.95" lane="1" heatid="21010" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="919" birthdate="2010-01-01" gender="F" lastname="Belger" firstname="Linnea" license="392772">
              <RESULTS>
                <RESULT resultid="4301" eventid="19" swimtime="00:00:51.02" lane="8" heatid="19018" />
                <RESULT resultid="4302" eventid="25" swimtime="00:00:47.96" lane="7" heatid="25010" />
                <RESULT resultid="4303" eventid="33" swimtime="00:01:27.18" lane="7" heatid="33006" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="920" birthdate="2014-01-01" gender="F" lastname="Grämer" firstname="Stella" license="445949">
              <RESULTS>
                <RESULT resultid="4304" eventid="17" swimtime="00:01:04.39" lane="5" heatid="17007" />
                <RESULT resultid="4305" eventid="21" swimtime="00:01:04.62" lane="6" heatid="21008" />
                <RESULT resultid="4306" eventid="25" swimtime="00:00:54.70" lane="5" heatid="25007" />
                <RESULT resultid="4307" eventid="29" swimtime="00:00:46.54" lane="6" heatid="29008" />
                <RESULT resultid="4308" eventid="31" swimtime="00:01:08.22" lane="2" heatid="31003" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="921" birthdate="2014-01-01" gender="F" lastname="Heinrich" firstname="Thea" license="445950">
              <RESULTS>
                <RESULT resultid="4309" eventid="19" swimtime="00:00:52.36" lane="6" heatid="19009" />
                <RESULT resultid="4310" eventid="25" swimtime="00:00:52.24" lane="6" heatid="25010" />
                <RESULT resultid="4311" eventid="27" swimtime="00:00:59.41" lane="1" heatid="27011" />
                <RESULT resultid="4312" eventid="29" swimtime="00:00:47.77" lane="2" heatid="29009" />
                <RESULT resultid="4313" eventid="33" swimtime="00:01:49.14" lane="2" heatid="33004" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="922" birthdate="2008-01-01" gender="M" lastname="Heinrich" firstname="Tim" license="364363">
              <RESULTS>
                <RESULT resultid="4314" eventid="4" swimtime="00:01:24.69" lane="4" heatid="4003" />
                <RESULT resultid="4315" eventid="6" swimtime="00:00:31.91" lane="1" heatid="6009" />
                <RESULT resultid="4316" eventid="13" swimtime="00:00:26.75" lane="3" heatid="13017" />
                <RESULT resultid="4317" eventid="20" swimtime="00:00:33.87" lane="5" heatid="20022" />
                <RESULT resultid="4318" eventid="26" swimtime="00:00:32.66" lane="7" heatid="26023" />
                <RESULT resultid="4319" eventid="34" swimtime="00:01:03.77" lane="2" heatid="34015" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="923" birthdate="2012-01-01" gender="F" lastname="Kaiser" firstname="Zoe" license="431997">
              <RESULTS>
                <RESULT resultid="4320" eventid="10" swimtime="00:01:41.00" lane="1" heatid="10006" />
                <RESULT resultid="4321" eventid="12" swimtime="00:00:36.53" lane="8" heatid="12009" />
                <RESULT resultid="4322" eventid="17" swimtime="00:00:50.75" lane="7" heatid="17016" />
                <RESULT resultid="4323" eventid="21" swimtime="00:00:51.14" lane="7" heatid="21014" />
                <RESULT resultid="4324" eventid="31" swimtime="00:00:55.03" lane="1" heatid="31006" />
                <RESULT resultid="4325" eventid="33" swimtime="00:01:20.62" lane="8" heatid="33008" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY number="1" gender="X" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="4234" eventid="7" swimtime="00:02:41.97" lane="1" heatid="7002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:28.00" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="923" number="1" />
                    <RELAYPOSITION athleteid="915" number="2" />
                    <RELAYPOSITION athleteid="906" number="3" />
                    <RELAYPOSITION athleteid="912" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB name="Dresdner Delphine e.V." nation="GER" region="12" code="5753">
          <ATHLETES>
            <ATHLETE athleteid="1157" birthdate="2010-01-01" gender="M" lastname="Dieckmann" firstname="Albert" license="409638">
              <RESULTS>
                <RESULT resultid="5423" eventid="2" swimtime="00:03:04.58" lane="2" heatid="2005">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:28.33" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="5424" eventid="11" swimtime="00:01:27.00" lane="5" heatid="11008" />
                <RESULT resultid="5425" eventid="13" swimtime="00:00:34.06" lane="7" heatid="13011" />
                <RESULT resultid="5426" eventid="20" swimtime="00:00:44.20" lane="6" heatid="20017" />
                <RESULT resultid="5427" eventid="26" swimtime="00:00:39.10" lane="7" heatid="26021" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1158" birthdate="2009-01-01" gender="M" lastname="Piotrowski" firstname="Alexej" license="467916">
              <RESULTS>
                <RESULT resultid="5428" eventid="6" swimtime="00:00:39.99" lane="4" heatid="6004" />
                <RESULT resultid="5429" eventid="13" status="DNS" swimtime="00:00:00.00" lane="8" heatid="13014" />
                <RESULT resultid="5430" eventid="34" swimtime="00:01:16.64" lane="8" heatid="34011" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1159" birthdate="2009-01-01" gender="F" lastname="Zubovska" firstname="Alina" license="454879">
              <RESULTS>
                <RESULT resultid="5431" eventid="5" swimtime="00:00:30.61" lane="6" heatid="5014" />
                <RESULT resultid="5432" eventid="12" swimtime="00:00:30.16" lane="3" heatid="12017" />
                <RESULT resultid="5433" eventid="23" swimtime="00:02:32.12" lane="5" heatid="23011">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:11.04" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="5434" eventid="33" swimtime="00:01:07.67" lane="1" heatid="33018" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1160" birthdate="2010-01-01" gender="F" lastname="Ratzenbeck" firstname="Amalia Maria" license="472042">
              <RESULTS>
                <RESULT resultid="5435" eventid="1" swimtime="00:02:54.56" lane="4" heatid="1006">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:25.63" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="5436" eventid="5" swimtime="00:00:35.10" lane="4" heatid="5012" />
                <RESULT resultid="5437" eventid="14" swimtime="00:03:11.45" lane="2" heatid="14007">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:32.96" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1161" birthdate="2013-01-01" gender="F" lastname="Henze" firstname="Anna" license="445341">
              <RESULTS>
                <RESULT resultid="5438" eventid="1" swimtime="00:03:24.19" lane="4" heatid="1002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:36.48" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="5439" eventid="5" swimtime="00:00:40.70" lane="5" heatid="5006" />
                <RESULT resultid="5440" eventid="10" swimtime="00:01:33.14" lane="4" heatid="10011" />
                <RESULT resultid="5441" eventid="12" swimtime="00:00:35.64" lane="7" heatid="12011" />
                <RESULT resultid="5442" eventid="17" swimtime="00:00:51.13" lane="1" heatid="17016" />
                <RESULT resultid="5443" eventid="25" swimtime="00:00:40.45" lane="6" heatid="25026" />
                <RESULT resultid="5444" eventid="31" swimtime="00:00:51.78" lane="7" heatid="31007" />
                <RESULT resultid="5445" eventid="37" swimtime="00:03:11.79" lane="1" heatid="37004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:36.25" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1162" birthdate="2014-01-01" gender="F" lastname="Pinera de la Cruz" firstname="Annika" license="447790">
              <RESULTS>
                <RESULT resultid="5446" eventid="17" swimtime="00:01:19.06" lane="3" heatid="17001" />
                <RESULT resultid="5447" eventid="19" swimtime="00:00:52.49" lane="1" heatid="19016" />
                <RESULT resultid="5448" eventid="25" swimtime="00:00:57.01" lane="2" heatid="25006" />
                <RESULT resultid="5449" eventid="27" swimtime="00:01:01.05" lane="3" heatid="27010" />
                <RESULT resultid="5450" eventid="29" swimtime="00:00:52.84" lane="3" heatid="29006" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1163" birthdate="2010-01-01" gender="M" lastname="Böhme" firstname="Anton" license="402826">
              <RESULTS>
                <RESULT resultid="5451" eventid="4" swimtime="00:01:24.71" lane="8" heatid="4011" />
                <RESULT resultid="5452" eventid="6" swimtime="00:00:36.92" lane="1" heatid="6008" />
                <RESULT resultid="5453" eventid="15" swimtime="00:02:56.64" lane="6" heatid="15007">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:26.49" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1164" birthdate="2009-01-01" gender="F" lastname="Rückert" firstname="Arja" license="395284">
              <RESULTS>
                <RESULT resultid="5454" eventid="5" swimtime="00:00:38.46" lane="5" heatid="5008" />
                <RESULT resultid="5455" eventid="10" swimtime="00:01:30.68" lane="2" heatid="10005" />
                <RESULT resultid="5456" eventid="12" swimtime="00:00:33.74" lane="8" heatid="12014" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1165" birthdate="2008-01-01" gender="M" lastname="Kessler" firstname="Arthur" license="448029">
              <RESULTS>
                <RESULT resultid="5457" eventid="6" status="DNS" swimtime="00:00:00.00" lane="6" heatid="6008" />
                <RESULT resultid="5458" eventid="13" status="DNS" swimtime="00:00:00.00" lane="8" heatid="13016" />
                <RESULT resultid="5459" eventid="34" status="DNS" swimtime="00:00:00.00" lane="2" heatid="34012" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1166" birthdate="2010-01-01" gender="F" lastname="Pinkert" firstname="Camilla" license="402824">
              <RESULTS>
                <RESULT resultid="5460" eventid="1" swimtime="00:03:12.98" lane="5" heatid="1002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:28.43" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="5461" eventid="5" swimtime="00:00:37.96" lane="5" heatid="5010" />
                <RESULT resultid="5462" eventid="12" swimtime="00:00:35.18" lane="2" heatid="12012" />
                <RESULT resultid="5463" eventid="23" swimtime="00:02:53.08" lane="1" heatid="23007">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:21.03" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1167" birthdate="2013-01-01" gender="F" lastname="Holstein" firstname="Carla" license="467930">
              <RESULTS>
                <RESULT resultid="5464" eventid="17" swimtime="00:01:19.16" lane="1" heatid="17003" />
                <RESULT resultid="5465" eventid="19" swimtime="00:00:57.24" lane="4" heatid="19009" />
                <RESULT resultid="5466" eventid="27" swimtime="00:01:08.06" lane="8" heatid="27001" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1168" birthdate="2014-01-01" gender="M" lastname="Hesse" firstname="Carlo" license="447796">
              <RESULTS>
                <RESULT resultid="5467" eventid="18" swimtime="00:01:01.32" lane="6" heatid="18009" />
                <RESULT resultid="5468" eventid="22" status="DSQ" swimtime="00:01:01.74" lane="8" heatid="22007" comment="Start vor dem Startsignal." />
                <RESULT resultid="5469" eventid="26" swimtime="00:00:50.56" lane="7" heatid="26008" />
                <RESULT resultid="5470" eventid="30" swimtime="00:00:54.69" lane="6" heatid="30003" />
                <RESULT resultid="5471" eventid="32" swimtime="00:01:12.59" lane="4" heatid="32001" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1169" birthdate="2013-01-01" gender="F" lastname="Grimm" firstname="Carmen" license="467466">
              <RESULTS>
                <RESULT resultid="5472" eventid="17" status="DNS" swimtime="00:00:00.00" lane="3" heatid="17002" />
                <RESULT resultid="5473" eventid="21" status="DNS" swimtime="00:00:00.00" lane="2" heatid="21007" />
                <RESULT resultid="5474" eventid="25" status="DNS" swimtime="00:00:00.00" lane="6" heatid="25012" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1170" birthdate="2013-01-01" gender="F" lastname="Böhmert" firstname="Charlotte Katrin" license="437495">
              <RESULTS>
                <RESULT resultid="5475" eventid="3" swimtime="00:01:54.66" lane="6" heatid="3004" />
                <RESULT resultid="5476" eventid="5" swimtime="00:00:46.17" lane="7" heatid="5004" />
                <RESULT resultid="5477" eventid="19" swimtime="00:00:51.61" lane="5" heatid="19017" />
                <RESULT resultid="5478" eventid="23" swimtime="00:03:25.54" lane="7" heatid="23002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:37.94" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="5479" eventid="33" swimtime="00:01:31.72" lane="4" heatid="33007" />
                <RESULT resultid="5480" eventid="37" swimtime="00:03:33.07" lane="6" heatid="37003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:44.20" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1171" birthdate="2014-01-01" gender="F" lastname="Ziller" firstname="Charlotte Wilhelmine" license="451281">
              <RESULTS>
                <RESULT resultid="5481" eventid="17" swimtime="00:01:03.40" lane="2" heatid="17014" />
                <RESULT resultid="5482" eventid="19" swimtime="00:00:56.01" lane="7" heatid="19011" />
                <RESULT resultid="5483" eventid="25" swimtime="00:00:48.53" lane="8" heatid="25020" />
                <RESULT resultid="5484" eventid="27" swimtime="00:01:04.33" lane="7" heatid="27003" />
                <RESULT resultid="5485" eventid="31" swimtime="00:01:05.61" lane="8" heatid="31005" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1172" birthdate="2006-01-01" gender="F" lastname="Römmermann" firstname="Chiara" license="348341">
              <RESULTS>
                <RESULT resultid="5486" eventid="5" swimtime="00:00:32.47" lane="1" heatid="5014" />
                <RESULT resultid="5487" eventid="10" swimtime="00:01:14.82" lane="7" heatid="10016" />
                <RESULT resultid="5488" eventid="23" swimtime="00:02:26.55" lane="7" heatid="23011">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:09.38" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="5489" eventid="33" swimtime="00:01:06.26" lane="5" heatid="33017" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1173" birthdate="2012-01-01" gender="F" lastname="Bambynek" firstname="Clara" license="437403">
              <RESULTS>
                <RESULT resultid="5490" eventid="3" swimtime="00:01:49.49" lane="2" heatid="3007" />
                <RESULT resultid="5491" eventid="10" swimtime="00:01:37.49" lane="8" heatid="10006" />
                <RESULT resultid="5492" eventid="14" swimtime="00:04:00.14" lane="1" heatid="14004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:55.97" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="5493" eventid="19" swimtime="00:00:46.51" lane="6" heatid="19022" />
                <RESULT resultid="5494" eventid="25" swimtime="00:00:44.65" lane="3" heatid="25021" />
                <RESULT resultid="5495" eventid="33" swimtime="00:01:29.76" lane="4" heatid="33006" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1174" birthdate="2009-01-01" gender="F" lastname="Gutberlet" firstname="Clara" license="395293">
              <RESULTS>
                <RESULT resultid="5496" eventid="1" swimtime="00:02:56.17" lane="7" heatid="1005">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:25.40" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="5497" eventid="14" swimtime="00:03:12.88" lane="8" heatid="14007">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:33.10" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="5498" eventid="19" swimtime="00:00:39.95" lane="6" heatid="19026" />
                <RESULT resultid="5499" eventid="23" swimtime="00:02:41.39" lane="4" heatid="23010">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:16.97" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1175" birthdate="2010-01-01" gender="F" lastname="Zimmerling" firstname="Clara" license="402811">
              <RESULTS>
                <RESULT resultid="5500" eventid="12" swimtime="00:00:28.04" lane="6" heatid="12018" />
                <RESULT resultid="5501" eventid="23" swimtime="00:02:17.18" lane="4" heatid="23011">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:03.84" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="5502" eventid="33" swimtime="00:01:02.08" lane="5" heatid="33018" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1176" birthdate="2011-01-01" gender="F" lastname="Dank" firstname="Daria" license="437415">
              <RESULTS>
                <RESULT resultid="5503" eventid="14" swimtime="00:03:57.99" lane="6" heatid="14002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:53.96" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="5504" eventid="19" swimtime="00:00:49.92" lane="4" heatid="19017" />
                <RESULT resultid="5505" eventid="25" swimtime="00:00:52.63" lane="3" heatid="25011" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1177" birthdate="2014-01-01" gender="F" lastname="Küllig" firstname="Ella Maria" license="449169">
              <RESULTS>
                <RESULT resultid="5506" eventid="17" swimtime="00:01:19.43" lane="3" heatid="17003" />
                <RESULT resultid="5507" eventid="19" swimtime="00:00:57.46" lane="2" heatid="19008" />
                <RESULT resultid="5508" eventid="25" swimtime="00:01:01.74" lane="7" heatid="25007" />
                <RESULT resultid="5509" eventid="27" swimtime="00:01:11.99" lane="8" heatid="27008" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1178" birthdate="2009-01-01" gender="M" lastname="Müller" firstname="Emil" license="395288">
              <RESULTS>
                <RESULT resultid="5510" eventid="24" swimtime="00:02:11.68" lane="5" heatid="24009">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:02.72" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="5511" eventid="34" swimtime="00:00:59.87" lane="6" heatid="34015" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1179" birthdate="2011-01-01" gender="M" lastname="Thätner" firstname="Erek" license="445404">
              <RESULTS>
                <RESULT resultid="5512" eventid="20" swimtime="00:00:49.32" lane="6" heatid="20012" />
                <RESULT resultid="5513" eventid="24" swimtime="00:03:11.57" lane="1" heatid="24003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:34.99" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="5514" eventid="26" swimtime="00:00:46.13" lane="1" heatid="26013" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1180" birthdate="2012-01-01" gender="M" lastname="Zimmerling" firstname="Erik" license="437405">
              <RESULTS>
                <RESULT resultid="5515" eventid="2" swimtime="00:02:59.27" lane="6" heatid="2006">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:26.16" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="5516" eventid="6" swimtime="00:00:38.27" lane="2" heatid="6007" />
                <RESULT resultid="5517" eventid="11" swimtime="00:01:21.36" lane="3" heatid="11010" />
                <RESULT resultid="5518" eventid="13" swimtime="00:00:31.95" lane="8" heatid="13013" />
                <RESULT resultid="5519" eventid="20" swimtime="00:00:40.74" lane="1" heatid="20020" />
                <RESULT resultid="5520" eventid="24" swimtime="00:02:47.13" lane="3" heatid="24007">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:19.82" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="5521" eventid="26" swimtime="00:00:35.59" lane="5" heatid="26022" />
                <RESULT resultid="5522" eventid="34" swimtime="00:01:12.14" lane="6" heatid="34012" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1181" birthdate="2012-01-01" gender="M" lastname="Krüger" firstname="Felix" license="437406">
              <RESULTS>
                <RESULT resultid="5523" eventid="4" swimtime="00:01:45.94" lane="2" heatid="4003" />
                <RESULT resultid="5524" eventid="11" swimtime="00:01:22.67" lane="6" heatid="11010" />
                <RESULT resultid="5525" eventid="13" swimtime="00:00:35.59" lane="7" heatid="13010" />
                <RESULT resultid="5526" eventid="15" swimtime="00:03:52.96" lane="4" heatid="15001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:52.52" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="5527" eventid="18" swimtime="00:00:50.38" lane="5" heatid="18012" />
                <RESULT resultid="5528" eventid="26" swimtime="00:00:38.39" lane="1" heatid="26022" />
                <RESULT resultid="5529" eventid="34" swimtime="00:01:22.16" lane="4" heatid="34009" />
                <RESULT resultid="5530" eventid="38" swimtime="00:02:56.05" lane="7" heatid="38004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:27.08" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1182" birthdate="2014-01-01" gender="F" lastname="Trodler" firstname="Felizia" license="447789">
              <RESULTS>
                <RESULT resultid="5531" eventid="17" swimtime="00:01:05.05" lane="8" heatid="17006" />
                <RESULT resultid="5532" eventid="19" swimtime="00:00:56.75" lane="7" heatid="19010" />
                <RESULT resultid="5533" eventid="25" swimtime="00:00:55.40" lane="3" heatid="25008" />
                <RESULT resultid="5534" eventid="27" swimtime="00:01:06.60" lane="2" heatid="27008" />
                <RESULT resultid="5535" eventid="29" swimtime="00:00:47.19" lane="7" heatid="29008" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1183" birthdate="2013-01-01" gender="M" lastname="Böhmert" firstname="Flinn Jan" license="437496">
              <RESULTS>
                <RESULT resultid="5536" eventid="2" swimtime="00:03:38.58" lane="7" heatid="2002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:44.56" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="5537" eventid="6" swimtime="00:00:48.10" lane="7" heatid="6002" />
                <RESULT resultid="5538" eventid="18" swimtime="00:00:53.55" lane="7" heatid="18012" />
                <RESULT resultid="5539" eventid="24" swimtime="00:03:17.82" lane="4" heatid="24002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:36.89" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="5540" eventid="34" swimtime="00:01:28.32" lane="1" heatid="34005" />
                <RESULT resultid="5541" eventid="38" swimtime="00:03:26.84" lane="4" heatid="38002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:42.35" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1184" birthdate="2013-01-01" gender="M" lastname="Köhler" firstname="Fritz" license="447788">
              <RESULTS>
                <RESULT resultid="5542" eventid="18" swimtime="00:01:09.73" lane="5" heatid="18006" />
                <RESULT resultid="5543" eventid="20" swimtime="00:00:59.36" lane="4" heatid="20004" />
                <RESULT resultid="5544" eventid="26" swimtime="00:00:57.30" lane="8" heatid="26006" />
                <RESULT resultid="5545" eventid="28" swimtime="00:01:10.00" lane="8" heatid="28004" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1185" birthdate="2012-01-01" gender="M" lastname="Hermann" firstname="Gregor" license="475074">
              <RESULTS>
                <RESULT resultid="5546" eventid="4" swimtime="00:02:03.65" lane="3" heatid="4001" />
                <RESULT resultid="5547" eventid="13" swimtime="00:00:49.17" lane="7" heatid="13001" />
                <RESULT resultid="5548" eventid="15" swimtime="00:04:24.92" lane="3" heatid="15001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:02:08.86" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1186" birthdate="2011-01-01" gender="F" lastname="Hollain" firstname="Greta" license="424864">
              <RESULTS>
                <RESULT resultid="5549" eventid="19" swimtime="00:00:46.49" lane="4" heatid="19016" />
                <RESULT resultid="5550" eventid="25" swimtime="00:00:46.09" lane="7" heatid="25019" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1187" birthdate="2014-01-01" gender="F" lastname="Böhmert" firstname="Hannah" license="447997">
              <RESULTS>
                <RESULT resultid="5551" eventid="17" swimtime="00:01:04.68" lane="7" heatid="17013" />
                <RESULT resultid="5552" eventid="19" swimtime="00:00:57.83" lane="3" heatid="19010" />
                <RESULT resultid="5553" eventid="25" swimtime="00:00:51.50" lane="6" heatid="25016" />
                <RESULT resultid="5554" eventid="29" swimtime="00:00:44.76" lane="4" heatid="29011" />
                <RESULT resultid="5555" eventid="31" swimtime="00:01:09.85" lane="3" heatid="31004" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1188" birthdate="2010-01-01" gender="F" lastname="Gärtner" firstname="Hannah" license="402813">
              <RESULTS>
                <RESULT resultid="5556" eventid="1" swimtime="00:03:08.38" lane="1" heatid="1005">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:28.22" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="5557" eventid="23" swimtime="00:02:49.48" lane="7" heatid="23009">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:18.00" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1189" birthdate="2014-01-01" gender="F" lastname="Krause" firstname="Helena" license="447793">
              <RESULTS>
                <RESULT resultid="5558" eventid="17" status="DSQ" swimtime="00:01:06.54" lane="1" heatid="17007" comment="Start vor dem Startsignal" />
                <RESULT resultid="5559" eventid="21" swimtime="00:00:59.11" lane="6" heatid="21010" />
                <RESULT resultid="5560" eventid="25" swimtime="00:00:53.04" lane="4" heatid="25011" />
                <RESULT resultid="5561" eventid="29" swimtime="00:00:44.48" lane="4" heatid="29010" />
                <RESULT resultid="5562" eventid="31" swimtime="00:01:12.34" lane="6" heatid="31003" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1190" birthdate="2007-01-01" gender="M" lastname="Sachs" firstname="Hermann" license="365266">
              <RESULTS>
                <RESULT resultid="5563" eventid="13" swimtime="00:00:28.74" lane="2" heatid="13016" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1191" birthdate="2012-01-01" gender="M" lastname="Jeschke" firstname="Jakob" license="437407">
              <RESULTS>
                <RESULT resultid="5564" eventid="2" swimtime="00:03:39.16" lane="2" heatid="2002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:43.14" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="5565" eventid="6" swimtime="00:00:45.40" lane="6" heatid="6003" />
                <RESULT resultid="5566" eventid="11" swimtime="00:01:43.73" lane="1" heatid="11004" />
                <RESULT resultid="5567" eventid="13" swimtime="00:00:38.54" lane="1" heatid="13004" />
                <RESULT resultid="5568" eventid="18" swimtime="00:00:58.93" lane="3" heatid="18010" />
                <RESULT resultid="5569" eventid="22" swimtime="00:00:55.70" lane="8" heatid="22009" />
                <RESULT resultid="5570" eventid="26" swimtime="00:00:44.51" lane="5" heatid="26013" />
                <RESULT resultid="5571" eventid="34" swimtime="00:01:29.58" lane="1" heatid="34004" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1192" birthdate="2013-01-01" gender="F" lastname="Hänig" firstname="Jasna" license="445403">
              <RESULTS>
                <RESULT resultid="5572" eventid="1" swimtime="00:03:25.92" lane="6" heatid="1003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:34.17" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="5573" eventid="5" swimtime="00:00:39.78" lane="2" heatid="5007" />
                <RESULT resultid="5574" eventid="10" swimtime="00:01:31.37" lane="8" heatid="10010" />
                <RESULT resultid="5575" eventid="12" swimtime="00:00:38.67" lane="3" heatid="12008" />
                <RESULT resultid="5576" eventid="21" swimtime="00:00:52.24" lane="5" heatid="21012" />
                <RESULT resultid="5577" eventid="23" swimtime="00:03:09.35" lane="7" heatid="23005">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:29.06" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="5578" eventid="33" swimtime="00:01:22.86" lane="6" heatid="33009" />
                <RESULT resultid="5579" eventid="37" status="DSQ" swimtime="00:03:21.78" lane="3" heatid="37001" comment="Bei der 3. Wende wurde die Wende nicht unverzüglich nach Einnahme der Bauchlage ausgeführt.">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:37.42" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1193" birthdate="2007-01-01" gender="M" lastname="Weigel" firstname="Joan-Maurice" license="365268">
              <RESULTS>
                <RESULT resultid="5580" eventid="4" swimtime="00:01:25.83" lane="5" heatid="4010" />
                <RESULT resultid="5581" eventid="13" swimtime="00:00:27.17" lane="4" heatid="13017" />
                <RESULT resultid="5582" eventid="20" swimtime="00:00:35.97" lane="4" heatid="20021" />
                <RESULT resultid="5583" eventid="34" swimtime="00:01:04.69" lane="3" heatid="34014" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1194" birthdate="2013-01-01" gender="M" lastname="Hänig" firstname="Johannes" license="437401">
              <RESULTS>
                <RESULT resultid="5584" eventid="4" swimtime="00:01:37.83" lane="1" heatid="4008" />
                <RESULT resultid="5585" eventid="11" swimtime="00:01:42.80" lane="5" heatid="11003" />
                <RESULT resultid="5586" eventid="13" swimtime="00:00:37.73" lane="6" heatid="13007" />
                <RESULT resultid="5587" eventid="15" swimtime="00:03:31.33" lane="1" heatid="15003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:44.12" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="5588" eventid="20" swimtime="00:00:43.11" lane="1" heatid="20018" />
                <RESULT resultid="5589" eventid="26" swimtime="00:00:45.85" lane="8" heatid="26015" />
                <RESULT resultid="5590" eventid="28" swimtime="00:00:51.27" lane="5" heatid="28008" />
                <RESULT resultid="5591" eventid="34" swimtime="00:01:29.48" lane="1" heatid="34007" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1195" birthdate="2011-01-01" gender="M" lastname="Schuricht" firstname="Jonas" license="473948">
              <RESULTS>
                <RESULT resultid="5592" eventid="13" status="DNS" swimtime="00:00:00.00" lane="6" heatid="13001" />
                <RESULT resultid="5593" eventid="26" swimtime="00:00:50.01" lane="4" heatid="26009" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1196" birthdate="2014-01-01" gender="F" lastname="Näther" firstname="Josephin" license="452213">
              <RESULTS>
                <RESULT resultid="5594" eventid="17" swimtime="00:00:59.91" lane="1" heatid="17008" />
                <RESULT resultid="5595" eventid="21" swimtime="00:01:00.09" lane="3" heatid="21006" />
                <RESULT resultid="5596" eventid="25" swimtime="00:00:50.29" lane="1" heatid="25013" />
                <RESULT resultid="5597" eventid="29" swimtime="00:00:48.29" lane="2" heatid="29006" />
                <RESULT resultid="5598" eventid="31" swimtime="00:01:11.29" lane="2" heatid="31002" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1197" birthdate="2014-01-01" gender="M" lastname="Walter" firstname="Julius" license="447798">
              <RESULTS>
                <RESULT resultid="5599" eventid="18" swimtime="00:00:54.44" lane="5" heatid="18011" />
                <RESULT resultid="5600" eventid="22" swimtime="00:00:53.40" lane="6" heatid="22009" />
                <RESULT resultid="5601" eventid="26" swimtime="00:00:47.94" lane="7" heatid="26011" />
                <RESULT resultid="5602" eventid="30" swimtime="00:00:46.75" lane="7" heatid="30006" />
                <RESULT resultid="5603" eventid="32" swimtime="00:01:05.19" lane="7" heatid="32003" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1198" birthdate="2011-01-01" gender="F" lastname="Wächter" firstname="Lara Helene" license="424860">
              <RESULTS>
                <RESULT resultid="5604" eventid="1" swimtime="00:03:40.80" lane="4" heatid="1001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:41.58" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="5605" eventid="5" swimtime="00:00:44.18" lane="4" heatid="5003" />
                <RESULT resultid="5606" eventid="12" swimtime="00:00:38.15" lane="3" heatid="12006" />
                <RESULT resultid="5607" eventid="25" swimtime="00:00:43.01" lane="7" heatid="25023" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1199" birthdate="2008-01-01" gender="F" lastname="Peter" firstname="Lara Marie" license="387128">
              <RESULTS>
                <RESULT resultid="5608" eventid="1" swimtime="00:02:59.11" lane="4" heatid="1005">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:23.66" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="5609" eventid="12" swimtime="00:00:31.60" lane="7" heatid="12017" />
                <RESULT resultid="5610" eventid="23" swimtime="00:02:34.65" lane="1" heatid="23011">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:13.57" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="5611" eventid="33" swimtime="00:01:11.34" lane="3" heatid="33017" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1200" birthdate="2012-01-01" gender="F" lastname="Drechsel" firstname="Lea Emilia" license="445397">
              <RESULTS>
                <RESULT resultid="5612" eventid="17" swimtime="00:01:03.99" lane="6" heatid="17009" />
                <RESULT resultid="5613" eventid="23" swimtime="00:03:15.66" lane="8" heatid="23002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:35.15" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="5614" eventid="33" swimtime="00:01:32.92" lane="2" heatid="33008" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1201" birthdate="2012-01-01" gender="F" lastname="Lähner" firstname="Lea" license="437408">
              <RESULTS>
                <RESULT resultid="5615" eventid="3" swimtime="00:01:57.37" lane="1" heatid="3004" />
                <RESULT resultid="5616" eventid="10" swimtime="00:01:52.96" lane="5" heatid="10002" />
                <RESULT resultid="5617" eventid="12" swimtime="00:00:42.82" lane="1" heatid="12004" />
                <RESULT resultid="5618" eventid="14" swimtime="00:04:05.58" lane="6" heatid="14001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:02:00.32" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="5619" eventid="19" swimtime="00:00:51.88" lane="8" heatid="19016" />
                <RESULT resultid="5620" eventid="21" swimtime="00:00:56.33" lane="2" heatid="21011" />
                <RESULT resultid="5621" eventid="25" swimtime="00:00:49.49" lane="8" heatid="25021" />
                <RESULT resultid="5622" eventid="33" swimtime="00:01:40.47" lane="6" heatid="33005" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1202" birthdate="2013-01-01" gender="M" lastname="Barthel" firstname="Lennard" license="437409">
              <RESULTS>
                <RESULT resultid="5623" eventid="2" swimtime="00:03:19.06" lane="3" heatid="2004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:34.60" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="5624" eventid="6" swimtime="00:00:39.47" lane="7" heatid="6006" />
                <RESULT resultid="5625" eventid="13" swimtime="00:00:35.01" lane="4" heatid="13007" />
                <RESULT resultid="5626" eventid="22" swimtime="00:00:51.11" lane="8" heatid="22011" />
                <RESULT resultid="5627" eventid="24" swimtime="00:03:00.66" lane="6" heatid="24005">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:27.60" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="5628" eventid="34" swimtime="00:01:21.18" lane="4" heatid="34008" />
                <RESULT resultid="5629" eventid="36" swimtime="00:01:37.27" lane="1" heatid="36002" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1203" birthdate="2014-01-01" gender="F" lastname="Jurke" firstname="Leonie Johanna" license="448038">
              <RESULTS>
                <RESULT resultid="5630" eventid="17" swimtime="00:01:13.46" lane="2" heatid="17002" />
                <RESULT resultid="5631" eventid="19" swimtime="00:00:51.48" lane="2" heatid="19014" />
                <RESULT resultid="5632" eventid="25" swimtime="00:00:49.16" lane="1" heatid="25009" />
                <RESULT resultid="5633" eventid="27" swimtime="00:00:58.14" lane="4" heatid="27010" />
                <RESULT resultid="5634" eventid="29" swimtime="00:00:45.61" lane="6" heatid="29009" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1204" birthdate="2012-01-01" gender="F" lastname="Sauer" firstname="Liesbeth" license="444965">
              <RESULTS>
                <RESULT resultid="5635" eventid="3" swimtime="00:01:33.30" lane="4" heatid="3009" />
                <RESULT resultid="6364" eventid="12" swimtime="00:00:33.34" lane="8" heatid="12002" />
                <RESULT resultid="5637" eventid="14" status="DNS" swimtime="00:00:00.00" lane="7" heatid="14006" />
                <RESULT resultid="5638" eventid="19" swimtime="00:00:42.28" lane="6" heatid="19024" />
                <RESULT resultid="6365" eventid="27" swimtime="00:00:52.05" lane="5" heatid="27002" />
                <RESULT resultid="5640" eventid="33" swimtime="00:01:14.94" lane="2" heatid="33015" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1205" birthdate="2012-01-01" gender="F" lastname="Vogel" firstname="Lina" license="437392">
              <RESULTS>
                <RESULT resultid="5642" eventid="3" swimtime="00:01:39.54" lane="3" heatid="3009" />
                <RESULT resultid="5643" eventid="10" swimtime="00:01:30.29" lane="1" heatid="10011" />
                <RESULT resultid="5644" eventid="14" swimtime="00:03:33.75" lane="6" heatid="14005">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:44.58" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="5645" eventid="19" swimtime="00:00:45.11" lane="1" heatid="19024" />
                <RESULT resultid="5646" eventid="25" swimtime="00:00:41.39" lane="1" heatid="25026" />
                <RESULT resultid="5647" eventid="33" swimtime="00:01:26.04" lane="5" heatid="33009" />
                <RESULT resultid="5648" eventid="37" swimtime="00:03:13.63" lane="4" heatid="37005">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:35.21" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1206" birthdate="2009-01-01" gender="F" lastname="Werner" firstname="Lotte" license="395286">
              <RESULTS>
                <RESULT resultid="5649" eventid="3" swimtime="00:01:34.76" lane="1" heatid="3010" />
                <RESULT resultid="5650" eventid="14" swimtime="00:03:21.87" lane="3" heatid="14006">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:37.21" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="5651" eventid="19" swimtime="00:00:42.27" lane="8" heatid="19026" />
                <RESULT resultid="5652" eventid="23" swimtime="00:02:47.91" lane="2" heatid="23009">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:19.06" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1207" birthdate="2015-01-01" gender="M" lastname="Egger" firstname="Luca" license="463555">
              <RESULTS>
                <RESULT resultid="5653" eventid="18" swimtime="00:01:00.32" lane="5" heatid="18010" />
                <RESULT resultid="5654" eventid="20" swimtime="00:00:57.39" lane="5" heatid="20008" />
                <RESULT resultid="5655" eventid="26" swimtime="00:00:48.37" lane="4" heatid="26012" />
                <RESULT resultid="5656" eventid="28" swimtime="00:01:05.48" lane="6" heatid="28006" />
                <RESULT resultid="5657" eventid="30" swimtime="00:00:45.35" lane="6" heatid="30007" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1208" birthdate="2010-01-01" gender="M" lastname="Schmidtke" firstname="Luca" license="402814">
              <RESULTS>
                <RESULT resultid="5658" eventid="2" swimtime="00:03:19.31" lane="1" heatid="2004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:34.57" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="5659" eventid="6" swimtime="00:00:41.37" lane="8" heatid="6006" />
                <RESULT resultid="5660" eventid="13" swimtime="00:00:33.89" lane="6" heatid="13011" />
                <RESULT resultid="5661" eventid="20" swimtime="00:00:46.46" lane="3" heatid="20013" />
                <RESULT resultid="5662" eventid="26" swimtime="00:00:41.33" lane="8" heatid="26020" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1209" birthdate="2009-01-01" gender="F" lastname="Liebs" firstname="Lucia Anita" license="395285">
              <RESULTS>
                <RESULT resultid="5663" eventid="1" swimtime="00:03:10.26" lane="5" heatid="1003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:33.15" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="5664" eventid="5" swimtime="00:00:38.37" lane="3" heatid="5009" />
                <RESULT resultid="5665" eventid="8" swimtime="00:03:32.09" lane="6" heatid="8001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:38.43" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="5666" eventid="25" swimtime="00:00:41.51" lane="7" heatid="25024" />
                <RESULT resultid="5667" eventid="35" swimtime="00:01:28.91" lane="4" heatid="35002" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1210" birthdate="2012-01-01" gender="F" lastname="Kovanovic" firstname="Maja" license="448554">
              <RESULTS>
                <RESULT resultid="5668" eventid="1" swimtime="00:03:27.79" lane="3" heatid="1002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:41.52" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="5669" eventid="3" swimtime="00:01:56.54" lane="7" heatid="3004" />
                <RESULT resultid="5670" eventid="10" swimtime="00:01:43.06" lane="5" heatid="10006" />
                <RESULT resultid="5671" eventid="14" swimtime="00:04:02.69" lane="1" heatid="14003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:57.41" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="5672" eventid="19" swimtime="00:00:53.83" lane="1" heatid="19017" />
                <RESULT resultid="5673" eventid="25" swimtime="00:00:45.34" lane="5" heatid="25022" />
                <RESULT resultid="5674" eventid="27" swimtime="00:01:02.62" lane="3" heatid="27009" />
                <RESULT resultid="5675" eventid="33" swimtime="00:01:31.64" lane="1" heatid="33008" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1211" birthdate="2014-01-01" gender="F" lastname="Richter" firstname="Marie-Sophie" license="446897">
              <RESULTS>
                <RESULT resultid="5676" eventid="19" swimtime="00:00:48.75" lane="5" heatid="19015" />
                <RESULT resultid="5677" eventid="21" swimtime="00:00:56.60" lane="8" heatid="21012" />
                <RESULT resultid="5678" eventid="25" swimtime="00:00:46.67" lane="1" heatid="25022" />
                <RESULT resultid="5679" eventid="29" swimtime="00:00:42.84" lane="6" heatid="29011" />
                <RESULT resultid="5680" eventid="31" swimtime="00:00:58.28" lane="5" heatid="31006" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1212" birthdate="2009-01-01" gender="M" lastname="Zielke" firstname="Mark Anthony" license="435533">
              <RESULTS>
                <RESULT resultid="5681" eventid="4" swimtime="00:01:36.27" lane="2" heatid="4008" />
                <RESULT resultid="5682" eventid="13" swimtime="00:00:33.68" lane="6" heatid="13010" />
                <RESULT resultid="5683" eventid="20" status="DNS" swimtime="00:00:00.00" lane="5" heatid="20019" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1213" birthdate="2012-01-01" gender="M" lastname="Haberkorn" firstname="Matthäus" license="437400">
              <RESULTS>
                <RESULT resultid="5684" eventid="2" swimtime="00:03:04.79" lane="7" heatid="2006">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:27.17" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="5685" eventid="6" swimtime="00:00:36.64" lane="4" heatid="6007" />
                <RESULT resultid="5686" eventid="11" swimtime="00:01:22.98" lane="2" heatid="11010" />
                <RESULT resultid="5687" eventid="13" swimtime="00:00:31.75" lane="3" heatid="13013" />
                <RESULT resultid="5688" eventid="20" status="DSQ" swimtime="00:00:44.61" lane="2" heatid="20014" comment="Mehrere Delphinkicks nach dem Start." />
                <RESULT resultid="5689" eventid="24" status="DSQ" swimtime="00:02:42.73" lane="6" heatid="24006" comment="Start vor dem Startsignal.">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:19.57" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="5690" eventid="26" swimtime="00:00:38.32" lane="7" heatid="26022" />
                <RESULT resultid="5691" eventid="34" swimtime="00:01:12.29" lane="7" heatid="34012" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1214" birthdate="2014-01-01" gender="M" lastname="Bambynek" firstname="Max" license="447791">
              <RESULTS>
                <RESULT resultid="5692" eventid="18" swimtime="00:01:04.60" lane="8" heatid="18008" />
                <RESULT resultid="5693" eventid="20" swimtime="00:00:55.72" lane="5" heatid="20007" />
                <RESULT resultid="5694" eventid="22" swimtime="00:01:03.31" lane="8" heatid="22006" />
                <RESULT resultid="5695" eventid="26" swimtime="00:00:49.80" lane="2" heatid="26011" />
                <RESULT resultid="5696" eventid="28" swimtime="00:01:04.89" lane="8" heatid="28006" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1215" birthdate="2011-01-01" gender="M" lastname="Gennerich" firstname="Maximilian" license="423096">
              <RESULTS>
                <RESULT resultid="5697" eventid="2" swimtime="00:02:43.10" lane="4" heatid="2007">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:20.42" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="5698" eventid="13" swimtime="00:00:29.87" lane="4" heatid="13014" />
                <RESULT resultid="5699" eventid="24" swimtime="00:02:23.94" lane="7" heatid="24009">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:09.40" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="5700" eventid="34" swimtime="00:01:05.33" lane="1" heatid="34014" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1216" birthdate="2008-01-01" gender="F" lastname="Kirsten" firstname="Melanie" license="406782">
              <RESULTS>
                <RESULT resultid="5701" eventid="10" status="WDR" swimtime="00:00:00.00" lane="7" heatid="10010" />
                <RESULT resultid="5702" eventid="12" status="WDR" swimtime="00:00:00.00" lane="7" heatid="12009" />
                <RESULT resultid="5703" eventid="25" status="WDR" swimtime="00:00:00.00" lane="4" heatid="25025" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1217" birthdate="2011-01-01" gender="F" lastname="Pöche" firstname="Mia" license="448550">
              <RESULTS>
                <RESULT resultid="5704" eventid="1" swimtime="00:03:39.44" lane="8" heatid="1002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:41.14" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="5705" eventid="5" swimtime="00:00:46.39" lane="8" heatid="5002" />
                <RESULT resultid="5706" eventid="12" swimtime="00:00:39.81" lane="7" heatid="12007" />
                <RESULT resultid="5707" eventid="23" swimtime="00:03:23.70" lane="2" heatid="23003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:35.00" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="5708" eventid="25" swimtime="00:00:45.29" lane="1" heatid="25023" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1218" birthdate="2012-01-01" gender="F" lastname="Müller" firstname="Milene" license="437414">
              <RESULTS>
                <RESULT resultid="5709" eventid="1" swimtime="00:03:05.81" lane="1" heatid="1006">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:26.49" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="5710" eventid="5" swimtime="00:00:36.65" lane="2" heatid="5010" />
                <RESULT resultid="5711" eventid="10" swimtime="00:01:23.40" lane="1" heatid="10014" />
                <RESULT resultid="5712" eventid="12" swimtime="00:00:32.38" lane="5" heatid="12014" />
                <RESULT resultid="5713" eventid="19" swimtime="00:00:42.62" lane="6" heatid="19025" />
                <RESULT resultid="5714" eventid="25" swimtime="00:00:37.81" lane="3" heatid="25033" />
                <RESULT resultid="5715" eventid="33" swimtime="00:01:14.23" lane="8" heatid="33016" />
                <RESULT resultid="5716" eventid="37" swimtime="00:02:57.04" lane="7" heatid="37007">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:27.34" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1219" birthdate="2012-01-01" gender="F" lastname="Neugebauer" firstname="Neele" license="448555">
              <RESULTS>
                <RESULT resultid="5717" eventid="3" swimtime="00:01:47.27" lane="6" heatid="3005" />
                <RESULT resultid="5718" eventid="5" swimtime="00:00:47.11" lane="2" heatid="5004" />
                <RESULT resultid="5719" eventid="10" swimtime="00:01:36.31" lane="1" heatid="10008" />
                <RESULT resultid="5720" eventid="14" swimtime="00:03:48.93" lane="5" heatid="14003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:52.89" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="5721" eventid="19" swimtime="00:00:47.95" lane="4" heatid="19018" />
                <RESULT resultid="5722" eventid="25" swimtime="00:00:41.85" lane="2" heatid="25023" />
                <RESULT resultid="5723" eventid="27" swimtime="00:01:00.13" lane="7" heatid="27010" />
                <RESULT resultid="5724" eventid="33" swimtime="00:01:26.13" lane="8" heatid="33010" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1220" birthdate="2013-01-01" gender="F" lastname="Engel" firstname="Nele Sunshine" license="466521">
              <RESULTS>
                <RESULT resultid="5725" eventid="17" swimtime="00:01:05.11" lane="6" heatid="17006" />
                <RESULT resultid="5726" eventid="19" swimtime="00:01:05.34" lane="1" heatid="19006" />
                <RESULT resultid="5727" eventid="21" swimtime="00:01:12.64" lane="7" heatid="21003" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1221" birthdate="2014-01-01" gender="M" lastname="Sonnabend" firstname="Nils" license="454545">
              <RESULTS>
                <RESULT resultid="5728" eventid="20" swimtime="00:00:52.58" lane="3" heatid="20009" />
                <RESULT resultid="5729" eventid="22" swimtime="00:00:50.24" lane="1" heatid="22011" />
                <RESULT resultid="5730" eventid="26" swimtime="00:00:47.70" lane="2" heatid="26012" />
                <RESULT resultid="5731" eventid="28" swimtime="00:01:01.27" lane="1" heatid="28006" />
                <RESULT resultid="5732" eventid="32" swimtime="00:00:56.64" lane="8" heatid="32005" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1222" birthdate="2009-01-01" gender="F" lastname="Bröse" firstname="Nora" license="395289">
              <RESULTS>
                <RESULT resultid="5733" eventid="10" swimtime="00:01:25.70" lane="2" heatid="10013" />
                <RESULT resultid="5734" eventid="12" swimtime="00:00:33.72" lane="3" heatid="12014" />
                <RESULT resultid="5735" eventid="23" swimtime="00:02:41.89" lane="6" heatid="23008">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:18.77" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="5736" eventid="25" swimtime="00:00:38.28" lane="2" heatid="25031" />
                <RESULT resultid="5737" eventid="33" swimtime="00:01:15.28" lane="7" heatid="33015" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1223" birthdate="2011-01-01" gender="M" lastname="Lieske" firstname="Oliver" license="424850">
              <RESULTS>
                <RESULT resultid="5738" eventid="2" swimtime="00:03:20.92" lane="1" heatid="2003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:33.55" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="5739" eventid="4" swimtime="00:01:46.64" lane="1" heatid="4006" />
                <RESULT resultid="5740" eventid="13" swimtime="00:00:36.10" lane="6" heatid="13009" />
                <RESULT resultid="5741" eventid="15" swimtime="00:03:54.95" lane="2" heatid="15004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:53.61" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1224" birthdate="2011-01-01" gender="M" lastname="Kurth" firstname="Otis" license="424846">
              <RESULTS>
                <RESULT resultid="5742" eventid="4" swimtime="00:01:38.45" lane="7" heatid="4007" />
                <RESULT resultid="5743" eventid="13" swimtime="00:00:31.36" lane="4" heatid="13012" />
                <RESULT resultid="5744" eventid="15" swimtime="00:03:37.17" lane="3" heatid="15004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:46.39" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1225" birthdate="2011-01-01" gender="M" lastname="Dieckmann" firstname="Patrick" license="424848">
              <RESULTS>
                <RESULT resultid="5745" eventid="2" swimtime="00:02:55.42" lane="5" heatid="2006">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:24.67" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="5746" eventid="6" swimtime="00:00:37.86" lane="6" heatid="6007" />
                <RESULT resultid="5747" eventid="11" swimtime="00:01:22.73" lane="7" heatid="11010" />
                <RESULT resultid="5748" eventid="13" swimtime="00:00:32.57" lane="6" heatid="13013" />
                <RESULT resultid="5749" eventid="20" swimtime="00:00:43.50" lane="3" heatid="20016" />
                <RESULT resultid="5750" eventid="24" swimtime="00:02:32.03" lane="6" heatid="24008">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:13.30" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="5751" eventid="26" swimtime="00:00:38.03" lane="5" heatid="26021" />
                <RESULT resultid="5752" eventid="38" swimtime="00:02:56.09" lane="6" heatid="38004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:24.43" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1226" birthdate="2014-01-01" gender="F" lastname="Haase" firstname="Paula" license="448182">
              <RESULTS>
                <RESULT resultid="5753" eventid="17" swimtime="00:01:07.74" lane="6" heatid="17005" />
                <RESULT resultid="5754" eventid="19" swimtime="00:00:55.86" lane="8" heatid="19011" />
                <RESULT resultid="5755" eventid="21" swimtime="00:01:00.26" lane="1" heatid="21009" />
                <RESULT resultid="5756" eventid="25" swimtime="00:00:54.20" lane="8" heatid="25012" />
                <RESULT resultid="5757" eventid="27" swimtime="00:01:02.49" lane="4" heatid="27008" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1227" birthdate="2011-01-01" gender="F" lastname="Thill" firstname="Paula" license="448547">
              <RESULTS>
                <RESULT resultid="5758" eventid="3" swimtime="00:01:45.16" lane="3" heatid="3007" />
                <RESULT resultid="5759" eventid="10" swimtime="00:01:34.65" lane="2" heatid="10006" />
                <RESULT resultid="5760" eventid="12" swimtime="00:00:39.09" lane="1" heatid="12005" />
                <RESULT resultid="5761" eventid="14" swimtime="00:03:57.34" lane="3" heatid="14003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:57.32" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="5762" eventid="19" swimtime="00:00:48.12" lane="8" heatid="19022" />
                <RESULT resultid="5763" eventid="25" swimtime="00:00:43.37" lane="4" heatid="25021" />
                <RESULT resultid="5764" eventid="33" swimtime="00:01:26.28" lane="4" heatid="33008" />
                <RESULT resultid="5765" eventid="37" swimtime="00:03:41.70" lane="5" heatid="37001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:50.93" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1228" birthdate="2008-01-01" gender="M" lastname="Meffert" firstname="Paule" license="379588">
              <RESULTS>
                <RESULT resultid="5766" eventid="13" swimtime="00:00:31.46" lane="3" heatid="13012" />
                <RESULT resultid="5767" eventid="15" swimtime="00:03:24.58" lane="4" heatid="15003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:31.80" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="5768" eventid="20" swimtime="00:00:37.63" lane="8" heatid="20021" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1229" birthdate="2013-01-01" gender="F" lastname="Balthasar" firstname="Paulina" license="452665">
              <RESULTS>
                <RESULT resultid="5769" eventid="12" status="DNS" swimtime="00:00:00.00" lane="6" heatid="12002" />
                <RESULT resultid="5770" eventid="17" swimtime="00:01:13.10" lane="6" heatid="17002" />
                <RESULT resultid="5771" eventid="21" swimtime="00:01:09.41" lane="1" heatid="21008" />
                <RESULT resultid="5772" eventid="25" swimtime="00:00:57.50" lane="8" heatid="25011" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1230" birthdate="2010-01-01" gender="F" lastname="Schreiber" firstname="Sarah" license="418099">
              <RESULTS>
                <RESULT resultid="5773" eventid="3" swimtime="00:01:38.85" lane="2" heatid="3008" />
                <RESULT resultid="5774" eventid="5" swimtime="00:00:44.45" lane="5" heatid="5005" />
                <RESULT resultid="5775" eventid="12" swimtime="00:00:38.79" lane="3" heatid="12007" />
                <RESULT resultid="5776" eventid="14" swimtime="00:03:36.38" lane="3" heatid="14005">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:44.99" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="5777" eventid="19" swimtime="00:00:45.31" lane="7" heatid="19022" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1231" birthdate="2013-01-01" gender="F" lastname="Lutcan" firstname="Stella" license="451942">
              <RESULTS>
                <RESULT resultid="5778" eventid="3" swimtime="00:02:09.95" lane="2" heatid="3002" />
                <RESULT resultid="5779" eventid="14" swimtime="00:04:28.04" lane="4" heatid="14001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:02:09.07" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="5780" eventid="17" swimtime="00:01:07.53" lane="4" heatid="17005" />
                <RESULT resultid="5781" eventid="19" swimtime="00:00:58.90" lane="2" heatid="19006" />
                <RESULT resultid="5782" eventid="25" swimtime="00:00:56.60" lane="8" heatid="25008" />
                <RESULT resultid="5783" eventid="27" swimtime="00:01:10.01" lane="1" heatid="27006" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1232" birthdate="2011-01-01" gender="F" lastname="Friese" firstname="Sunna Björk" license="448552">
              <RESULTS>
                <RESULT resultid="5784" eventid="3" swimtime="00:01:50.39" lane="5" heatid="3003" />
                <RESULT resultid="5785" eventid="5" swimtime="00:00:50.40" lane="6" heatid="5003" />
                <RESULT resultid="5786" eventid="12" swimtime="00:00:38.07" lane="6" heatid="12006" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1233" birthdate="2011-01-01" gender="F" lastname="Trodler" firstname="Tamara" license="424858">
              <RESULTS>
                <RESULT resultid="5787" eventid="3" swimtime="00:01:43.35" lane="4" heatid="3007" />
                <RESULT resultid="5788" eventid="10" swimtime="00:01:30.55" lane="2" heatid="10009" />
                <RESULT resultid="5789" eventid="12" swimtime="00:00:34.51" lane="3" heatid="12012" />
                <RESULT resultid="5790" eventid="19" swimtime="00:00:46.56" lane="3" heatid="19020" />
                <RESULT resultid="5791" eventid="23" swimtime="00:02:53.51" lane="6" heatid="23007">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:23.99" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="5792" eventid="33" swimtime="00:01:17.52" lane="6" heatid="33012" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1234" birthdate="2012-01-01" gender="F" lastname="Stillfried" firstname="Tara" license="437395">
              <RESULTS>
                <RESULT resultid="5793" eventid="5" swimtime="00:00:51.22" lane="2" heatid="5002" />
                <RESULT resultid="5794" eventid="10" swimtime="00:01:46.32" lane="6" heatid="10002" />
                <RESULT resultid="5795" eventid="12" swimtime="00:00:41.63" lane="4" heatid="12002" />
                <RESULT resultid="5796" eventid="25" swimtime="00:00:48.10" lane="2" heatid="25017" />
                <RESULT resultid="5797" eventid="27" swimtime="00:01:07.26" lane="4" heatid="27007" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1235" birthdate="2010-01-01" gender="F" lastname="Bil" firstname="Tjara Charleen" license="402823">
              <RESULTS>
                <RESULT resultid="5798" eventid="1" swimtime="00:03:04.70" lane="5" heatid="1005">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:22.20" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="5799" eventid="5" swimtime="00:00:33.86" lane="2" heatid="5013" />
                <RESULT resultid="5800" eventid="12" swimtime="00:00:32.52" lane="2" heatid="12016" />
                <RESULT resultid="5801" eventid="23" swimtime="00:02:43.51" lane="2" heatid="23006">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:18.07" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1236" birthdate="2012-01-01" gender="M" lastname="Sparka" firstname="Tom David" license="437398">
              <RESULTS>
                <RESULT resultid="5802" eventid="11" swimtime="00:01:33.46" lane="3" heatid="11006" />
                <RESULT resultid="5803" eventid="13" swimtime="00:00:38.61" lane="4" heatid="13005" />
                <RESULT resultid="5804" eventid="18" swimtime="00:00:55.30" lane="8" heatid="18011" />
                <RESULT resultid="5805" eventid="20" swimtime="00:00:50.42" lane="7" heatid="20010" />
                <RESULT resultid="5806" eventid="26" swimtime="00:00:43.12" lane="5" heatid="26017" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1237" birthdate="2012-01-01" gender="M" lastname="Örmeci" firstname="Ulas Kutay" license="448546">
              <RESULTS>
                <RESULT resultid="5807" eventid="4" swimtime="00:02:07.75" lane="7" heatid="4002" />
                <RESULT resultid="5808" eventid="13" swimtime="00:00:52.78" lane="2" heatid="13001" />
                <RESULT resultid="5809" eventid="15" swimtime="00:04:36.45" lane="7" heatid="15002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:02:16.12" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="5810" eventid="18" swimtime="00:01:27.98" lane="3" heatid="18002" />
                <RESULT resultid="5811" eventid="20" swimtime="00:00:58.36" lane="4" heatid="20005" />
                <RESULT resultid="5812" eventid="26" swimtime="00:00:58.67" lane="1" heatid="26004" />
                <RESULT resultid="5813" eventid="28" swimtime="00:01:05.70" lane="8" heatid="28003" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1238" birthdate="2012-01-01" gender="M" lastname="Ratzenbeck" firstname="Wilhelm David" license="472041">
              <RESULTS>
                <RESULT resultid="5814" eventid="2" swimtime="00:02:58.94" lane="8" heatid="2006">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:28.84" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="5815" eventid="4" swimtime="00:01:29.73" lane="7" heatid="4009" />
                <RESULT resultid="5816" eventid="15" swimtime="00:03:18.42" lane="3" heatid="15005">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:38.55" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1239" birthdate="2012-01-01" gender="F" lastname="Dong" firstname="Xichen" license="475075">
              <RESULTS>
                <RESULT resultid="5817" eventid="17" swimtime="00:01:13.05" lane="2" heatid="17001" />
                <RESULT resultid="5818" eventid="21" swimtime="00:01:03.75" lane="8" heatid="21002" />
                <RESULT resultid="5819" eventid="25" swimtime="00:00:56.03" lane="4" heatid="25001" />
                <RESULT resultid="5820" eventid="33" swimtime="00:02:07.57" lane="3" heatid="33001" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY number="1" gender="X" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="5419" eventid="16" swimtime="00:02:05.67" lane="6" heatid="16002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:07.17" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1190" number="1" />
                    <RELAYPOSITION athleteid="1193" number="2" />
                    <RELAYPOSITION athleteid="1159" number="3" />
                    <RELAYPOSITION athleteid="1178" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" gender="X" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="5420" eventid="7" swimtime="00:02:22.49" lane="3" heatid="7003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:16.26" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1180" number="1" />
                    <RELAYPOSITION athleteid="1163" number="2" />
                    <RELAYPOSITION athleteid="1160" number="3" />
                    <RELAYPOSITION athleteid="1235" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="2" gender="X" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="5421" eventid="16" swimtime="00:02:26.73" lane="5" heatid="16001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:16.58" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1222" number="1" />
                    <RELAYPOSITION athleteid="1228" number="2" />
                    <RELAYPOSITION athleteid="1209" number="3" />
                    <RELAYPOSITION athleteid="1199" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="2" gender="X" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="5422" eventid="7" swimtime="00:02:39.23" lane="3" heatid="7002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:25.85" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1233" number="1" />
                    <RELAYPOSITION athleteid="1230" number="2" />
                    <RELAYPOSITION athleteid="1208" number="3" />
                    <RELAYPOSITION athleteid="1224" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB name="Dresdner SC 1898" nation="GER" region="12" code="3332">
          <ATHLETES>
            <ATHLETE athleteid="1246" birthdate="2013-01-01" gender="F" lastname="Heinze" firstname="Abigail Louise" license="443667">
              <RESULTS>
                <RESULT resultid="5827" eventid="3" swimtime="00:01:53.41" lane="1" heatid="3005" />
                <RESULT resultid="5828" eventid="10" status="DSQ" swimtime="00:01:46.81" lane="4" heatid="10004" comment="Nach verlassen der Rückenlage Wende nicht unverzüglich eingeleitet." />
                <RESULT resultid="5829" eventid="12" swimtime="00:00:41.97" lane="4" heatid="12005" />
                <RESULT resultid="5830" eventid="14" swimtime="00:03:47.45" lane="5" heatid="14002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:50.90" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="5831" eventid="19" swimtime="00:00:49.91" lane="5" heatid="19016" />
                <RESULT resultid="5832" eventid="27" swimtime="00:00:54.13" lane="5" heatid="27011" />
                <RESULT resultid="5833" eventid="33" swimtime="00:01:30.73" lane="1" heatid="33006" />
                <RESULT resultid="5834" eventid="37" status="DSQ" swimtime="00:03:39.81" lane="4" heatid="37001" comment="Bei der 1. Wende wurde die Wende nicht unverzüglich nach Einnahme der Bauchlage ausgeführt.">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:52.44" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1247" birthdate="2008-01-01" gender="M" lastname="Zische" firstname="Adrian" license="380817">
              <RESULTS>
                <RESULT resultid="5835" eventid="4" swimtime="00:01:09.62" lane="4" heatid="4011" />
                <RESULT resultid="5836" eventid="15" swimtime="00:02:36.63" lane="4" heatid="15007">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:14.68" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1248" birthdate="2013-01-01" gender="M" lastname="Niekisch" firstname="Alexander" license="443679">
              <RESULTS>
                <RESULT resultid="5837" eventid="18" swimtime="00:00:56.53" lane="2" heatid="18011" />
                <RESULT resultid="5838" eventid="26" swimtime="00:00:42.20" lane="5" heatid="26016" />
                <RESULT resultid="5839" eventid="34" swimtime="00:01:24.34" lane="5" heatid="34004" />
                <RESULT resultid="5840" eventid="36" swimtime="00:01:45.84" lane="5" heatid="36001" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1249" birthdate="2012-01-01" gender="F" lastname="Kirberger" firstname="Alexandra" license="436906">
              <RESULTS>
                <RESULT resultid="5841" eventid="5" swimtime="00:00:36.50" lane="4" heatid="5008" />
                <RESULT resultid="5842" eventid="10" swimtime="00:01:26.47" lane="6" heatid="10012" />
                <RESULT resultid="5843" eventid="12" swimtime="00:00:37.51" lane="1" heatid="12007" />
                <RESULT resultid="5844" eventid="23" swimtime="00:02:51.64" lane="4" heatid="23006">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:23.89" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="5845" eventid="25" swimtime="00:00:40.70" lane="6" heatid="25024" />
                <RESULT resultid="5846" eventid="31" swimtime="00:00:52.46" lane="2" heatid="31007" />
                <RESULT resultid="5847" eventid="37" swimtime="00:02:59.75" lane="8" heatid="37006">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:29.13" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1250" birthdate="2012-01-01" gender="M" lastname="Chaplygin" firstname="Alexej" license="443662">
              <RESULTS>
                <RESULT resultid="5848" eventid="4" swimtime="00:01:57.64" lane="1" heatid="4002" />
                <RESULT resultid="5849" eventid="11" swimtime="00:01:36.33" lane="2" heatid="11004" />
                <RESULT resultid="5850" eventid="13" swimtime="00:00:41.89" lane="4" heatid="13002" />
                <RESULT resultid="5851" eventid="18" swimtime="00:00:51.27" lane="2" heatid="18012" />
                <RESULT resultid="5852" eventid="22" swimtime="00:00:52.52" lane="4" heatid="22010" />
                <RESULT resultid="5853" eventid="26" swimtime="00:00:44.35" lane="5" heatid="26012" />
                <RESULT resultid="5854" eventid="34" swimtime="00:01:32.07" lane="7" heatid="34002" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1251" birthdate="2015-01-01" gender="F" lastname="Schreck" firstname="Alma" license="463729">
              <RESULTS>
                <RESULT resultid="5855" eventid="17" swimtime="00:01:28.64" lane="6" heatid="17001" />
                <RESULT resultid="5856" eventid="19" swimtime="00:01:03.24" lane="6" heatid="19001" />
                <RESULT resultid="5857" eventid="25" swimtime="00:01:01.75" lane="1" heatid="25007" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1252" birthdate="2012-01-01" gender="F" lastname="Schwamberger" firstname="Alma" license="443041">
              <RESULTS>
                <RESULT resultid="5858" eventid="17" swimtime="00:01:14.26" lane="5" heatid="17004" />
                <RESULT resultid="5859" eventid="19" swimtime="00:00:50.40" lane="4" heatid="19013" />
                <RESULT resultid="5860" eventid="25" swimtime="00:00:51.17" lane="2" heatid="25018" />
                <RESULT resultid="5861" eventid="27" swimtime="00:01:00.02" lane="4" heatid="27009" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1253" birthdate="2014-01-01" gender="F" lastname="Schmelter" firstname="Alwine" license="463385">
              <RESULTS>
                <RESULT resultid="5862" eventid="17" swimtime="00:01:07.20" lane="5" heatid="17010" />
                <RESULT resultid="5863" eventid="25" swimtime="00:00:55.07" lane="6" heatid="25013" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1254" birthdate="2014-01-01" gender="F" lastname="Gutjahr" firstname="Anna Lena" license="448021">
              <RESULTS>
                <RESULT resultid="5864" eventid="19" swimtime="00:00:56.50" lane="5" heatid="19010" />
                <RESULT resultid="5865" eventid="21" swimtime="00:00:55.86" lane="1" heatid="21011" />
                <RESULT resultid="5866" eventid="25" swimtime="00:00:44.27" lane="5" heatid="25018" />
                <RESULT resultid="5867" eventid="29" swimtime="00:00:39.79" lane="4" heatid="29012" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1255" birthdate="2014-01-01" gender="F" lastname="Mathiszik" firstname="Anna" license="448117">
              <RESULTS>
                <RESULT resultid="5868" eventid="19" swimtime="00:00:58.82" lane="6" heatid="19005" />
                <RESULT resultid="5869" eventid="25" swimtime="00:00:57.44" lane="6" heatid="25008" />
                <RESULT resultid="5870" eventid="27" swimtime="00:01:12.03" lane="7" heatid="27005" />
                <RESULT resultid="5871" eventid="29" swimtime="00:00:56.35" lane="6" heatid="29003" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1256" birthdate="2009-01-01" gender="F" lastname="Wagenknecht" firstname="Anne- Felicia" license="395546">
              <RESULTS>
                <RESULT resultid="5872" eventid="1" swimtime="00:03:01.61" lane="6" heatid="1005">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:23.67" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="5873" eventid="5" swimtime="00:00:36.66" lane="7" heatid="5010" />
                <RESULT resultid="5874" eventid="12" swimtime="00:00:33.06" lane="4" heatid="12015" />
                <RESULT resultid="5875" eventid="23" swimtime="00:02:46.73" lane="1" heatid="23009">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:17.61" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="5876" eventid="33" swimtime="00:01:12.99" lane="4" heatid="33015" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1257" birthdate="2009-01-01" gender="F" lastname="Zische" firstname="Annika" license="393879">
              <RESULTS>
                <RESULT resultid="5877" eventid="14" swimtime="00:02:43.89" lane="4" heatid="14007">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:18.84" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="5878" eventid="35" swimtime="00:01:09.65" lane="4" heatid="35004" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1258" birthdate="2010-01-01" gender="M" lastname="Hanke" firstname="Arthur" license="444305">
              <RESULTS>
                <RESULT resultid="5879" eventid="2" swimtime="00:03:15.05" lane="3" heatid="2005">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:31.16" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="5880" eventid="4" swimtime="00:01:41.64" lane="3" heatid="4007" />
                <RESULT resultid="5881" eventid="11" swimtime="00:01:30.43" lane="5" heatid="11007" />
                <RESULT resultid="5882" eventid="13" swimtime="00:00:36.03" lane="7" heatid="13009" />
                <RESULT resultid="5883" eventid="20" swimtime="00:00:44.17" lane="6" heatid="20015" />
                <RESULT resultid="5884" eventid="26" swimtime="00:00:40.10" lane="2" heatid="26018" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1259" birthdate="2013-01-01" gender="M" lastname="Lange" firstname="Arthur" license="443672">
              <RESULTS>
                <RESULT resultid="5885" eventid="2" swimtime="00:03:28.50" lane="4" heatid="2002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:36.91" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="5886" eventid="6" swimtime="00:00:40.49" lane="6" heatid="6004" />
                <RESULT resultid="5887" eventid="11" swimtime="00:01:34.90" lane="6" heatid="11006" />
                <RESULT resultid="5888" eventid="13" swimtime="00:00:39.00" lane="2" heatid="13004" />
                <RESULT resultid="5889" eventid="18" swimtime="00:00:53.32" lane="3" heatid="18011" />
                <RESULT resultid="5890" eventid="22" swimtime="00:00:56.03" lane="1" heatid="22009" />
                <RESULT resultid="5891" eventid="26" swimtime="00:00:41.68" lane="1" heatid="26018" />
                <RESULT resultid="5892" eventid="34" swimtime="00:01:29.02" lane="5" heatid="34003" />
                <RESULT resultid="5893" eventid="38" swimtime="00:03:17.47" lane="5" heatid="38002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:37.54" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1260" birthdate="2010-01-01" gender="M" lastname="Draganov" firstname="Atanas" license="427768">
              <RESULTS>
                <RESULT resultid="5894" eventid="2" swimtime="00:03:34.04" lane="3" heatid="2002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:38.95" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="5895" eventid="4" swimtime="00:01:58.00" lane="4" heatid="4002" />
                <RESULT resultid="5896" eventid="6" swimtime="00:00:44.35" lane="3" heatid="6004" />
                <RESULT resultid="5897" eventid="13" swimtime="00:00:35.86" lane="2" heatid="13007" />
                <RESULT resultid="5898" eventid="24" swimtime="00:03:10.61" lane="7" heatid="24003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:29.60" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="5899" eventid="26" swimtime="00:00:42.01" lane="7" heatid="26018" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1261" birthdate="2009-01-01" gender="M" lastname="Wüstenhagen" firstname="Aurel" license="395576">
              <RESULTS>
                <RESULT resultid="5900" eventid="2" swimtime="00:02:27.67" lane="5" heatid="2008">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:08.29" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="5901" eventid="13" swimtime="00:00:27.69" lane="2" heatid="13017" />
                <RESULT resultid="5902" eventid="24" swimtime="00:02:08.36" lane="3" heatid="24009">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:01.06" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="5903" eventid="34" swimtime="00:00:59.99" lane="3" heatid="34015" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1262" birthdate="2014-01-01" gender="M" lastname="Salfitzky" firstname="Benno" license="448061">
              <RESULTS>
                <RESULT resultid="5904" eventid="18" swimtime="00:00:54.19" lane="8" heatid="18012" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1263" birthdate="2014-01-01" gender="F" lastname="Harnisch" firstname="Carlotta" license="448039">
              <RESULTS>
                <RESULT resultid="5905" eventid="17" swimtime="00:00:59.53" lane="4" heatid="17009" />
                <RESULT resultid="5906" eventid="21" swimtime="00:01:01.76" lane="2" heatid="21008" />
                <RESULT resultid="5907" eventid="25" swimtime="00:00:44.66" lane="1" heatid="25021" />
                <RESULT resultid="5908" eventid="29" swimtime="00:00:44.63" lane="4" heatid="29009" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1264" birthdate="2015-01-01" gender="F" lastname="Matthes" firstname="Charlotte" license="463217">
              <RESULTS>
                <RESULT resultid="5909" eventid="17" status="WDR" swimtime="00:00:00.00" lane="8" heatid="17013" />
                <RESULT resultid="5910" eventid="19" status="WDR" swimtime="00:00:00.00" lane="8" heatid="19005" />
                <RESULT resultid="5911" eventid="25" status="WDR" swimtime="00:00:00.00" lane="4" heatid="25015" />
                <RESULT resultid="5912" eventid="29" status="WDR" swimtime="00:00:00.00" lane="3" heatid="29008" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1265" birthdate="2009-01-01" gender="F" lastname="Streiber" firstname="Charlotte" license="398189">
              <RESULTS>
                <RESULT resultid="5913" eventid="5" swimtime="00:00:34.83" lane="3" heatid="5011" />
                <RESULT resultid="5914" eventid="12" swimtime="00:00:32.56" lane="8" heatid="12016" />
                <RESULT resultid="5915" eventid="23" swimtime="00:02:38.24" lane="5" heatid="23009">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:16.24" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="5916" eventid="33" swimtime="00:01:12.13" lane="2" heatid="33016" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1266" birthdate="2009-01-01" gender="F" lastname="von Bonin" firstname="Charlotte" license="393877">
              <RESULTS>
                <RESULT resultid="5917" eventid="3" swimtime="00:01:35.71" lane="5" heatid="3008" />
                <RESULT resultid="5918" eventid="5" swimtime="00:00:37.55" lane="7" heatid="5009" />
                <RESULT resultid="5919" eventid="10" swimtime="00:01:24.48" lane="5" heatid="10010" />
                <RESULT resultid="5920" eventid="12" swimtime="00:00:33.99" lane="5" heatid="12013" />
                <RESULT resultid="5921" eventid="19" swimtime="00:00:44.28" lane="1" heatid="19023" />
                <RESULT resultid="5922" eventid="25" swimtime="00:00:38.87" lane="5" heatid="25027" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1267" birthdate="2010-01-01" gender="M" lastname="Schubert" firstname="Christian" license="412734">
              <RESULTS>
                <RESULT resultid="5923" eventid="2" swimtime="00:02:30.43" lane="3" heatid="2008">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:12.00" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="5924" eventid="6" swimtime="00:00:33.56" lane="2" heatid="6009" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1268" birthdate="2013-01-01" gender="F" lastname="Rotzsch" firstname="Clara Paulina" license="448155">
              <RESULTS>
                <RESULT resultid="5925" eventid="17" swimtime="00:00:59.50" lane="5" heatid="17008" />
                <RESULT resultid="5926" eventid="19" swimtime="00:00:55.64" lane="2" heatid="19015" />
                <RESULT resultid="5927" eventid="23" swimtime="00:03:46.40" lane="5" heatid="23001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:47.09" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="5928" eventid="27" swimtime="00:01:12.13" lane="2" heatid="27004" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1269" birthdate="2012-01-01" gender="F" lastname="Seidel" firstname="Dana" license="436901">
              <RESULTS>
                <RESULT resultid="5929" eventid="3" swimtime="00:01:46.51" lane="3" heatid="3005" />
                <RESULT resultid="5930" eventid="5" swimtime="00:00:44.12" lane="8" heatid="5005" />
                <RESULT resultid="5931" eventid="10" swimtime="00:01:31.74" lane="2" heatid="10010" />
                <RESULT resultid="5932" eventid="12" swimtime="00:00:36.86" lane="5" heatid="12008" />
                <RESULT resultid="5933" eventid="21" swimtime="00:00:52.53" lane="2" heatid="21014" />
                <RESULT resultid="5934" eventid="23" swimtime="00:03:02.33" lane="4" heatid="23005">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:28.88" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="5935" eventid="35" swimtime="00:01:47.00" lane="1" heatid="35002" />
                <RESULT resultid="5936" eventid="37" swimtime="00:03:18.94" lane="2" heatid="37003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:39.72" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1270" birthdate="2012-01-01" gender="M" lastname="Kolkowski" firstname="Daniel" license="443040">
              <RESULTS>
                <RESULT resultid="5937" eventid="2" swimtime="00:03:17.30" lane="7" heatid="2004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:31.21" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="5938" eventid="6" swimtime="00:00:40.55" lane="6" heatid="6005" />
                <RESULT resultid="5939" eventid="11" swimtime="00:01:25.53" lane="8" heatid="11009" />
                <RESULT resultid="5940" eventid="13" swimtime="00:00:36.50" lane="4" heatid="13009" />
                <RESULT resultid="5941" eventid="24" swimtime="00:02:50.21" lane="1" heatid="24007">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:21.05" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="5942" eventid="26" swimtime="00:00:39.23" lane="3" heatid="26019" />
                <RESULT resultid="5943" eventid="34" swimtime="00:01:18.58" lane="3" heatid="34010" />
                <RESULT resultid="5944" eventid="38" swimtime="00:02:54.44" lane="1" heatid="38004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:27.39" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1271" birthdate="2013-01-01" gender="M" lastname="Ulbricht" firstname="Daniel" license="443686">
              <RESULTS>
                <RESULT resultid="5945" eventid="20" swimtime="00:00:49.81" lane="8" heatid="20011" />
                <RESULT resultid="5946" eventid="24" swimtime="00:03:06.35" lane="1" heatid="24005">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:27.84" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="5947" eventid="32" swimtime="00:01:05.03" lane="8" heatid="32003" />
                <RESULT resultid="5948" eventid="38" swimtime="00:03:12.70" lane="3" heatid="38002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:34.09" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1272" birthdate="2013-01-01" gender="M" lastname="Khavrus" firstname="Dmitri" license="443668">
              <RESULTS>
                <RESULT resultid="5949" eventid="2" swimtime="00:03:23.69" lane="6" heatid="2003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:41.98" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="5950" eventid="4" swimtime="00:01:40.82" lane="3" heatid="4006" />
                <RESULT resultid="5951" eventid="13" swimtime="00:00:35.60" lane="6" heatid="13008" />
                <RESULT resultid="5952" eventid="15" swimtime="00:03:44.01" lane="1" heatid="15004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:49.77" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="5953" eventid="20" swimtime="00:00:44.34" lane="4" heatid="20014" />
                <RESULT resultid="5954" eventid="26" swimtime="00:00:40.29" lane="7" heatid="26019" />
                <RESULT resultid="5955" eventid="34" swimtime="00:01:18.28" lane="6" heatid="34007" />
                <RESULT resultid="5956" eventid="38" swimtime="00:03:14.21" lane="4" heatid="38001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:36.45" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1273" birthdate="2014-01-01" gender="M" lastname="Granzow" firstname="Edward" license="448232">
              <RESULTS>
                <RESULT resultid="5957" eventid="18" swimtime="00:01:06.14" lane="4" heatid="18005" />
                <RESULT resultid="5958" eventid="22" swimtime="00:01:08.75" lane="8" heatid="22004" />
                <RESULT resultid="5959" eventid="28" swimtime="00:01:20.34" lane="8" heatid="28002" />
                <RESULT resultid="5960" eventid="30" swimtime="00:00:46.79" lane="4" heatid="30004" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1274" birthdate="2009-01-01" gender="F" lastname="Packenius" firstname="Elena" license="396078">
              <RESULTS>
                <RESULT resultid="5961" eventid="1" swimtime="00:02:56.18" lane="7" heatid="1006">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:21.22" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="5962" eventid="5" swimtime="00:00:35.24" lane="2" heatid="5011" />
                <RESULT resultid="5963" eventid="19" swimtime="00:00:43.17" lane="5" heatid="19024" />
                <RESULT resultid="5964" eventid="33" swimtime="00:01:12.57" lane="6" heatid="33014" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1275" birthdate="2015-01-01" gender="F" lastname="Kirchner" firstname="Ella" license="463200">
              <RESULTS>
                <RESULT resultid="5965" eventid="17" swimtime="00:00:59.88" lane="3" heatid="17015" />
                <RESULT resultid="5966" eventid="19" swimtime="00:00:52.60" lane="7" heatid="19004" />
                <RESULT resultid="5967" eventid="25" swimtime="00:00:45.37" lane="4" heatid="25020" />
                <RESULT resultid="5968" eventid="29" swimtime="00:00:44.58" lane="1" heatid="29011" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1276" birthdate="2015-01-01" gender="M" lastname="Lieske" firstname="Emil" license="463225">
              <RESULTS>
                <RESULT resultid="5969" eventid="18" swimtime="00:01:14.24" lane="5" heatid="18003" />
                <RESULT resultid="5970" eventid="20" swimtime="00:01:19.40" lane="7" heatid="20001" />
                <RESULT resultid="5971" eventid="26" swimtime="00:01:03.41" lane="4" heatid="26002" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1277" birthdate="2012-01-01" gender="F" lastname="Stange" firstname="Emilia" license="436920">
              <RESULTS>
                <RESULT resultid="5972" eventid="5" swimtime="00:00:46.88" lane="3" heatid="5003" />
                <RESULT resultid="5973" eventid="10" swimtime="00:01:38.27" lane="3" heatid="10008" />
                <RESULT resultid="5974" eventid="17" swimtime="00:01:01.97" lane="1" heatid="17011" />
                <RESULT resultid="5975" eventid="25" swimtime="00:00:43.20" lane="6" heatid="25023" />
                <RESULT resultid="5976" eventid="33" swimtime="00:01:31.65" lane="6" heatid="33006" />
                <RESULT resultid="5977" eventid="37" status="DSQ" swimtime="00:03:23.21" lane="8" heatid="37003" comment="Bei der 3. Wende wurde die Wende nicht unverzüglich nach Einnahme der Bauchlage ausgeführt.">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:38.00" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1278" birthdate="2011-01-01" gender="M" lastname="Di Vincenzo" firstname="Emilio" license="436898">
              <RESULTS>
                <RESULT resultid="5978" eventid="20" status="WDR" swimtime="00:00:00.00" lane="1" heatid="20007" />
                <RESULT resultid="5979" eventid="26" status="WDR" swimtime="00:00:00.00" lane="5" heatid="26010" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1279" birthdate="2015-01-01" gender="F" lastname="Uebel" firstname="Emily" license="463205">
              <RESULTS>
                <RESULT resultid="5980" eventid="19" swimtime="00:01:00.81" lane="4" heatid="19004" />
                <RESULT resultid="5981" eventid="21" swimtime="00:01:03.71" lane="2" heatid="21009" />
                <RESULT resultid="5982" eventid="25" swimtime="00:00:56.14" lane="5" heatid="25010" />
                <RESULT resultid="5983" eventid="29" swimtime="00:00:52.56" lane="8" heatid="29005" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1280" birthdate="2015-01-01" gender="M" lastname="Böhme" firstname="Endrik" license="463193">
              <RESULTS>
                <RESULT resultid="5984" eventid="20" swimtime="00:01:07.90" lane="4" heatid="20002" />
                <RESULT resultid="5985" eventid="26" swimtime="00:01:04.15" lane="5" heatid="26002" />
                <RESULT resultid="5986" eventid="28" swimtime="00:01:10.91" lane="6" heatid="28002" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1281" birthdate="2015-01-01" gender="M" lastname="Beckmann" firstname="Erik" license="463196">
              <RESULTS>
                <RESULT resultid="5987" eventid="18" swimtime="00:01:16.15" lane="7" heatid="18004" />
                <RESULT resultid="5988" eventid="22" swimtime="00:01:17.44" lane="6" heatid="22004" />
                <RESULT resultid="5989" eventid="26" swimtime="00:00:58.43" lane="8" heatid="26004" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1282" birthdate="2015-01-01" gender="M" lastname="Schellhammer" firstname="Fabian" license="463209">
              <RESULTS>
                <RESULT resultid="5990" eventid="18" swimtime="00:01:09.04" lane="5" heatid="18007" />
                <RESULT resultid="5991" eventid="20" swimtime="00:01:07.00" lane="8" heatid="20001" />
                <RESULT resultid="5992" eventid="22" swimtime="00:01:13.31" lane="2" heatid="22005" />
                <RESULT resultid="5993" eventid="26" swimtime="00:01:01.90" lane="7" heatid="26005" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1283" birthdate="2014-01-01" gender="M" lastname="Kluge" firstname="Felix" license="449664">
              <RESULTS>
                <RESULT resultid="5994" eventid="18" swimtime="00:01:03.49" lane="7" heatid="18006" />
                <RESULT resultid="5995" eventid="20" swimtime="00:00:58.92" lane="8" heatid="20006" />
                <RESULT resultid="5996" eventid="22" swimtime="00:01:05.76" lane="5" heatid="22004" />
                <RESULT resultid="5997" eventid="28" swimtime="00:01:06.58" lane="7" heatid="28004" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1284" birthdate="2009-01-01" gender="M" lastname="Mehner" firstname="Felix" license="395569">
              <RESULTS>
                <RESULT resultid="5998" eventid="6" swimtime="00:00:32.24" lane="1" heatid="6010" />
                <RESULT resultid="5999" eventid="13" swimtime="00:00:28.24" lane="8" heatid="13017" />
                <RESULT resultid="6000" eventid="26" swimtime="00:00:32.08" lane="6" heatid="26024" />
                <RESULT resultid="6001" eventid="34" swimtime="00:01:03.42" lane="5" heatid="34014" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1285" birthdate="2011-01-01" gender="F" lastname="Auerswald" firstname="Florentine" license="424902">
              <RESULTS>
                <RESULT resultid="6002" eventid="3" swimtime="00:01:45.61" lane="8" heatid="3006" />
                <RESULT resultid="6003" eventid="5" swimtime="00:00:54.63" lane="4" heatid="5001" />
                <RESULT resultid="6004" eventid="12" swimtime="00:00:50.63" lane="5" heatid="12001" />
                <RESULT resultid="6005" eventid="14" swimtime="00:03:44.31" lane="2" heatid="14002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:48.09" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1286" birthdate="2015-01-01" gender="F" lastname="Kirberger" firstname="Franziska" license="463223">
              <RESULTS>
                <RESULT resultid="6006" eventid="17" swimtime="00:01:03.24" lane="3" heatid="17012" />
                <RESULT resultid="6007" eventid="19" swimtime="00:00:58.98" lane="8" heatid="19007" />
                <RESULT resultid="6008" eventid="21" swimtime="00:01:06.95" lane="7" heatid="21007" />
                <RESULT resultid="6009" eventid="27" swimtime="00:01:12.49" lane="1" heatid="27005" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1287" birthdate="2012-01-01" gender="M" lastname="Schiller" firstname="Fredo Matheo" license="436894">
              <RESULTS>
                <RESULT resultid="6010" eventid="20" swimtime="00:00:50.09" lane="7" heatid="20011" />
                <RESULT resultid="6011" eventid="28" swimtime="00:00:59.96" lane="7" heatid="28007" />
                <RESULT resultid="6012" eventid="32" swimtime="00:00:58.35" lane="7" heatid="32005" />
                <RESULT resultid="6013" eventid="34" swimtime="00:01:32.03" lane="8" heatid="34005" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1288" birthdate="2015-01-01" gender="M" lastname="Deichmüller" firstname="Friedrich" license="463211">
              <RESULTS>
                <RESULT resultid="6014" eventid="18" swimtime="00:01:09.34" lane="6" heatid="18006" />
                <RESULT resultid="6015" eventid="22" swimtime="00:01:08.45" lane="5" heatid="22003" />
                <RESULT resultid="6016" eventid="26" swimtime="00:00:55.11" lane="2" heatid="26006" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1289" birthdate="2008-01-01" gender="M" lastname="Drzymala" firstname="Fynn Mario" license="380796">
              <RESULTS>
                <RESULT resultid="6017" eventid="6" swimtime="00:00:26.90" lane="4" heatid="6011" />
                <RESULT resultid="6018" eventid="13" swimtime="00:00:26.37" lane="2" heatid="13018" />
                <RESULT resultid="6019" eventid="24" swimtime="00:02:05.19" lane="4" heatid="24009">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:58.83" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="6020" eventid="36" swimtime="00:01:00.00" lane="4" heatid="36003" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1290" birthdate="2012-01-01" gender="F" lastname="Sachse" firstname="Greta" license="436912">
              <RESULTS>
                <RESULT resultid="6021" eventid="3" swimtime="00:01:48.94" lane="4" heatid="3005" />
                <RESULT resultid="6022" eventid="5" swimtime="00:00:56.42" lane="1" heatid="5003" />
                <RESULT resultid="6023" eventid="12" swimtime="00:00:41.72" lane="7" heatid="12005" />
                <RESULT resultid="6024" eventid="14" swimtime="00:03:42.41" lane="4" heatid="14003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:50.18" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="6025" eventid="19" swimtime="00:00:47.26" lane="8" heatid="19019" />
                <RESULT resultid="6026" eventid="21" swimtime="00:00:58.95" lane="5" heatid="21009" />
                <RESULT resultid="6027" eventid="27" swimtime="00:00:56.20" lane="4" heatid="27011" />
                <RESULT resultid="6028" eventid="35" swimtime="00:02:07.64" lane="3" heatid="35001" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1291" birthdate="2011-01-01" gender="M" lastname="Winkler" firstname="Hannes" license="424910">
              <RESULTS>
                <RESULT resultid="6029" eventid="4" swimtime="00:01:48.54" lane="7" heatid="4004" />
                <RESULT resultid="6030" eventid="6" status="DSQ" swimtime="00:00:48.82" lane="8" heatid="6002" comment="Brustbeinbewegungen während der gesamten Schwimmstrecke." />
                <RESULT resultid="6031" eventid="11" swimtime="00:01:49.84" lane="4" heatid="11001" />
                <RESULT resultid="6032" eventid="13" swimtime="00:00:43.06" lane="2" heatid="13002" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1292" birthdate="2012-01-01" gender="F" lastname="Hanel" firstname="Heidi" license="436913">
              <RESULTS>
                <RESULT resultid="6033" eventid="1" swimtime="00:03:22.40" lane="1" heatid="1003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:31.05" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="6034" eventid="5" swimtime="00:00:39.53" lane="4" heatid="5005" />
                <RESULT resultid="6035" eventid="10" swimtime="00:01:26.78" lane="8" heatid="10013" />
                <RESULT resultid="6036" eventid="12" swimtime="00:00:34.70" lane="7" heatid="12012" />
                <RESULT resultid="6037" eventid="17" swimtime="00:00:48.08" lane="3" heatid="17016" />
                <RESULT resultid="6038" eventid="25" swimtime="00:00:37.84" lane="2" heatid="25032" />
                <RESULT resultid="6039" eventid="33" swimtime="00:01:24.12" lane="4" heatid="33009" />
                <RESULT resultid="6040" eventid="37" swimtime="00:03:07.99" lane="2" heatid="37005">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:33.46" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1293" birthdate="2008-01-01" gender="F" lastname="Göde" firstname="Helena" license="391855">
              <RESULTS>
                <RESULT resultid="6041" eventid="5" swimtime="00:00:28.82" lane="4" heatid="5014" />
                <RESULT resultid="6042" eventid="12" swimtime="00:00:27.96" lane="5" heatid="12018" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1294" birthdate="2013-01-01" gender="F" lastname="Hartmann" firstname="Helena" license="448024">
              <RESULTS>
                <RESULT resultid="6043" eventid="17" swimtime="00:01:03.21" lane="7" heatid="17008" />
                <RESULT resultid="6044" eventid="21" swimtime="00:01:02.55" lane="6" heatid="21004" />
                <RESULT resultid="6045" eventid="23" swimtime="00:03:50.48" lane="3" heatid="23001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:49.76" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="6046" eventid="27" swimtime="00:01:25.86" lane="6" heatid="27002" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1295" birthdate="2013-01-01" gender="F" lastname="Ragotzki" firstname="Helena" license="443681">
              <RESULTS>
                <RESULT resultid="6047" eventid="3" swimtime="00:01:57.12" lane="6" heatid="3002" />
                <RESULT resultid="6048" eventid="10" swimtime="00:01:48.87" lane="7" heatid="10004" />
                <RESULT resultid="6049" eventid="12" swimtime="00:00:43.76" lane="2" heatid="12003" />
                <RESULT resultid="6050" eventid="17" swimtime="00:00:56.56" lane="1" heatid="17014" />
                <RESULT resultid="6051" eventid="21" swimtime="00:00:56.85" lane="1" heatid="21012" />
                <RESULT resultid="6052" eventid="25" swimtime="00:00:49.21" lane="3" heatid="25016" />
                <RESULT resultid="6053" eventid="37" swimtime="00:03:44.78" lane="6" heatid="37001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:50.56" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1296" birthdate="2014-01-01" gender="F" lastname="Starke" firstname="Helene" license="449687">
              <RESULTS>
                <RESULT resultid="6054" eventid="17" swimtime="00:01:05.23" lane="8" heatid="17001" />
                <RESULT resultid="6055" eventid="19" swimtime="00:00:53.43" lane="3" heatid="19008" />
                <RESULT resultid="6056" eventid="25" swimtime="00:00:51.54" lane="4" heatid="25008" />
                <RESULT resultid="6057" eventid="29" swimtime="00:00:51.66" lane="4" heatid="29004" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1297" birthdate="2014-01-01" gender="F" lastname="Fischer" firstname="Henriette" license="448040">
              <RESULTS>
                <RESULT resultid="6058" eventid="17" swimtime="00:01:01.59" lane="8" heatid="17012" />
                <RESULT resultid="6059" eventid="21" swimtime="00:01:02.44" lane="4" heatid="21010" />
                <RESULT resultid="6060" eventid="25" swimtime="00:00:46.42" lane="1" heatid="25017" />
                <RESULT resultid="6061" eventid="29" swimtime="00:00:45.90" lane="2" heatid="29010" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1298" birthdate="2012-01-01" gender="F" lastname="Kobus" firstname="Henrijette" license="439567">
              <RESULTS>
                <RESULT resultid="6062" eventid="1" swimtime="00:02:45.18" lane="6" heatid="1007">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:16.99" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="6063" eventid="5" swimtime="00:00:32.92" lane="8" heatid="5014" />
                <RESULT resultid="6064" eventid="10" swimtime="00:01:16.21" lane="3" heatid="10015" />
                <RESULT resultid="6065" eventid="12" swimtime="00:00:30.13" lane="4" heatid="12017" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1299" birthdate="2015-01-01" gender="M" lastname="Schöbel" firstname="Jaden Dean" license="463206">
              <RESULTS>
                <RESULT resultid="6066" eventid="18" swimtime="00:01:14.55" lane="3" heatid="18006" />
                <RESULT resultid="6067" eventid="20" swimtime="00:01:05.89" lane="6" heatid="20002" />
                <RESULT resultid="6068" eventid="26" swimtime="00:01:02.95" lane="6" heatid="26003" />
                <RESULT resultid="6069" eventid="28" swimtime="00:01:12.19" lane="1" heatid="28003" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1300" birthdate="2013-01-01" gender="F" lastname="Suha" firstname="Jasmin" license="443682">
              <RESULTS>
                <RESULT resultid="6070" eventid="17" status="DSQ" swimtime="00:00:55.71" lane="4" heatid="17014" comment="Die wurden beim Anschlag nicht übereinander gehalten." />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1301" birthdate="2015-01-01" gender="M" lastname="Reichel" firstname="Johann Frederik" license="463208">
              <RESULTS>
                <RESULT resultid="6071" eventid="20" swimtime="00:01:04.33" lane="4" heatid="20001" />
                <RESULT resultid="6072" eventid="28" swimtime="00:01:11.81" lane="4" heatid="28003" />
                <RESULT resultid="6073" eventid="30" swimtime="00:01:02.68" lane="2" heatid="30001" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1302" birthdate="2015-01-01" gender="F" lastname="Obst" firstname="Johanna" license="463473">
              <RESULTS>
                <RESULT resultid="6074" eventid="17" swimtime="00:01:17.08" lane="1" heatid="17004" />
                <RESULT resultid="6075" eventid="21" swimtime="00:01:19.89" lane="3" heatid="21003" />
                <RESULT resultid="6076" eventid="25" swimtime="00:00:58.21" lane="1" heatid="25005" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1303" birthdate="2011-01-01" gender="F" lastname="Sachse" firstname="Johanna" license="424894">
              <RESULTS>
                <RESULT resultid="6077" eventid="3" swimtime="00:01:58.63" lane="1" heatid="3003" />
                <RESULT resultid="6078" eventid="10" swimtime="00:01:45.49" lane="1" heatid="10005" />
                <RESULT resultid="6079" eventid="12" swimtime="00:00:45.19" lane="1" heatid="12003" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1304" birthdate="2008-01-01" gender="M" lastname="Schmitt" firstname="Johannes" license="443043">
              <RESULTS>
                <RESULT resultid="6080" eventid="4" swimtime="00:01:29.98" lane="1" heatid="4010" />
                <RESULT resultid="6081" eventid="13" swimtime="00:00:30.58" lane="8" heatid="13015" />
                <RESULT resultid="6082" eventid="20" swimtime="00:00:38.74" lane="4" heatid="20020" />
                <RESULT resultid="6083" eventid="26" swimtime="00:00:39.12" lane="2" heatid="26020" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1305" birthdate="2014-01-01" gender="F" lastname="Barthel-Krauße" firstname="Jolien" license="463382">
              <RESULTS>
                <RESULT resultid="6084" eventid="17" swimtime="00:01:10.01" lane="3" heatid="17008" />
                <RESULT resultid="6085" eventid="19" swimtime="00:01:13.17" lane="2" heatid="19002" />
                <RESULT resultid="6086" eventid="29" swimtime="00:00:52.87" lane="6" heatid="29004" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1306" birthdate="2015-01-01" gender="F" lastname="Haas" firstname="Jolien" license="465085">
              <RESULTS>
                <RESULT resultid="6087" eventid="19" status="WDR" swimtime="00:00:00.00" lane="8" heatid="19003" />
                <RESULT resultid="6088" eventid="25" status="WDR" swimtime="00:00:00.00" lane="1" heatid="25004" />
                <RESULT resultid="6089" eventid="27" status="WDR" swimtime="00:00:00.00" lane="5" heatid="27000" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1307" birthdate="2015-01-01" gender="F" lastname="Hartmann" firstname="Josefine" license="463210">
              <RESULTS>
                <RESULT resultid="6090" eventid="19" swimtime="00:01:09.48" lane="6" heatid="19002" />
                <RESULT resultid="6091" eventid="25" swimtime="00:00:59.32" lane="6" heatid="25005" />
                <RESULT resultid="6092" eventid="27" status="DSQ" swimtime="00:01:23.65" lane="1" heatid="27001" comment="Das Brett wurde beim Zielsanschlag nicht vollständig umfasst." />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1308" birthdate="2014-01-01" gender="F" lastname="Schabel" firstname="Josefine" license="463198">
              <RESULTS>
                <RESULT resultid="6093" eventid="17" swimtime="00:01:19.21" lane="5" heatid="17003" />
                <RESULT resultid="6094" eventid="19" swimtime="00:01:10.66" lane="8" heatid="19004" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1309" birthdate="2009-01-01" gender="M" lastname="Lutter" firstname="Justus" license="419190">
              <RESULTS>
                <RESULT resultid="6095" eventid="6" swimtime="00:00:35.33" lane="3" heatid="6007" />
                <RESULT resultid="6096" eventid="13" swimtime="00:00:31.74" lane="1" heatid="13012" />
                <RESULT resultid="6097" eventid="20" swimtime="00:00:41.79" lane="3" heatid="20017" />
                <RESULT resultid="6098" eventid="34" swimtime="00:01:13.55" lane="7" heatid="34010" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1310" birthdate="2012-01-01" gender="M" lastname="Fritzsche" firstname="Karl" license="445371">
              <RESULTS>
                <RESULT resultid="6099" eventid="4" swimtime="00:01:44.31" lane="6" heatid="4005" />
                <RESULT resultid="6100" eventid="11" swimtime="00:01:44.76" lane="3" heatid="11002" />
                <RESULT resultid="6101" eventid="13" swimtime="00:00:43.28" lane="1" heatid="13003" />
                <RESULT resultid="6102" eventid="15" swimtime="00:03:54.08" lane="4" heatid="15002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:55.96" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1311" birthdate="2015-01-01" gender="M" lastname="Lages" firstname="Karl Hugo" license="463216">
              <RESULTS>
                <RESULT resultid="6103" eventid="18" swimtime="00:01:04.90" lane="2" heatid="18008" />
                <RESULT resultid="6104" eventid="20" status="DSQ" swimtime="00:01:01.98" lane="7" heatid="20002" comment="2 Delphinkicks" />
                <RESULT resultid="6105" eventid="26" swimtime="00:00:55.83" lane="4" heatid="26005" />
                <RESULT resultid="6106" eventid="30" swimtime="00:00:58.24" lane="3" heatid="30002" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1312" birthdate="2013-01-01" gender="F" lastname="Franke" firstname="Kim Sophie" license="443664">
              <RESULTS>
                <RESULT resultid="6107" eventid="17" swimtime="00:00:52.77" lane="5" heatid="17015" />
                <RESULT resultid="6108" eventid="25" swimtime="00:00:42.01" lane="8" heatid="25025" />
                <RESULT resultid="6109" eventid="33" swimtime="00:01:25.13" lane="3" heatid="33008" />
                <RESULT resultid="6110" eventid="37" swimtime="00:03:19.47" lane="4" heatid="37004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:37.72" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1313" birthdate="2015-01-01" gender="F" lastname="Beckmann" firstname="Klara" license="463195">
              <RESULTS>
                <RESULT resultid="6111" eventid="19" swimtime="00:01:00.94" lane="2" heatid="19005" />
                <RESULT resultid="6112" eventid="25" swimtime="00:00:59.57" lane="3" heatid="25006" />
                <RESULT resultid="6113" eventid="29" swimtime="00:00:59.04" lane="3" heatid="29003" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1314" birthdate="2010-01-01" gender="F" lastname="Dunkel" firstname="Lena" license="410626">
              <RESULTS>
                <RESULT resultid="6114" eventid="10" swimtime="00:01:15.85" lane="4" heatid="10015" />
                <RESULT resultid="6115" eventid="33" swimtime="00:01:10.54" lane="3" heatid="33016" />
                <RESULT resultid="6116" eventid="37" swimtime="00:02:43.41" lane="3" heatid="37007">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:20.15" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1315" birthdate="2010-01-01" gender="M" lastname="Martin" firstname="Levi" license="424888">
              <RESULTS>
                <RESULT resultid="6117" eventid="4" status="WDR" swimtime="00:00:00.00" lane="8" heatid="4008" />
                <RESULT resultid="6118" eventid="6" status="WDR" swimtime="00:00:00.00" lane="7" heatid="6003" />
                <RESULT resultid="6119" eventid="13" status="WDR" swimtime="00:00:00.00" lane="5" heatid="13006" />
                <RESULT resultid="6120" eventid="20" status="WDR" swimtime="00:00:00.00" lane="4" heatid="20015" />
                <RESULT resultid="6121" eventid="26" status="WDR" swimtime="00:00:00.00" lane="7" heatid="26013" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1316" birthdate="2015-01-01" gender="M" lastname="Otti" firstname="Lino" license="464258">
              <RESULTS>
                <RESULT resultid="6122" eventid="20" swimtime="00:01:00.87" lane="6" heatid="20005" />
                <RESULT resultid="6123" eventid="28" swimtime="00:01:14.09" lane="7" heatid="28003" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1317" birthdate="2013-01-01" gender="M" lastname="Wolf" firstname="Lio Maximilian" license="443688">
              <RESULTS>
                <RESULT resultid="6124" eventid="4" swimtime="00:01:59.75" lane="8" heatid="4003" />
                <RESULT resultid="6125" eventid="6" swimtime="00:00:57.22" lane="3" heatid="6001" />
                <RESULT resultid="6126" eventid="11" status="DSQ" swimtime="00:01:43.64" lane="7" heatid="11003" comment="Der Sportler leitete nach Verlassen der Rückenlage nicht unverzüglich die Wende ein." />
                <RESULT resultid="6127" eventid="13" swimtime="00:00:41.19" lane="8" heatid="13004" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1318" birthdate="2015-01-01" gender="F" lastname="Brüll" firstname="Lydia" license="463215">
              <RESULTS>
                <RESULT resultid="6128" eventid="17" swimtime="00:01:03.59" lane="7" heatid="17007" />
                <RESULT resultid="6129" eventid="21" swimtime="00:01:02.55" lane="8" heatid="21011" />
                <RESULT resultid="6130" eventid="25" swimtime="00:01:02.05" lane="8" heatid="25006" />
                <RESULT resultid="6131" eventid="27" status="DSQ" swimtime="00:01:22.05" lane="3" heatid="27002" comment="Wechselbeinschläge nach dem Start." />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1319" birthdate="2015-01-01" gender="F" lastname="Martin" firstname="Lykka-Marie" license="463227">
              <RESULTS>
                <RESULT resultid="6132" eventid="17" swimtime="00:01:16.04" lane="2" heatid="17004" />
                <RESULT resultid="6133" eventid="19" swimtime="00:01:06.84" lane="1" heatid="19002" />
                <RESULT resultid="6134" eventid="25" swimtime="00:01:02.15" lane="7" heatid="25004" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1320" birthdate="2011-01-01" gender="F" lastname="Winkler" firstname="Maike" license="424911">
              <RESULTS>
                <RESULT resultid="6135" eventid="1" swimtime="00:02:35.73" lane="3" heatid="1007">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:13.11" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="6136" eventid="5" swimtime="00:00:30.98" lane="2" heatid="5014" />
                <RESULT resultid="6137" eventid="12" swimtime="00:00:29.86" lane="1" heatid="12018" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1321" birthdate="2009-01-01" gender="F" lastname="Dörfer" firstname="Maja" license="393881">
              <RESULTS>
                <RESULT resultid="6138" eventid="1" swimtime="00:03:03.66" lane="3" heatid="1005">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:23.99" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="6139" eventid="5" swimtime="00:00:34.01" lane="6" heatid="5012" />
                <RESULT resultid="6140" eventid="25" swimtime="00:00:34.84" lane="2" heatid="25034" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1322" birthdate="2009-01-01" gender="M" lastname="Pöschmann" firstname="Marec" license="415182">
              <RESULTS>
                <RESULT resultid="6141" eventid="13" swimtime="00:00:27.89" lane="8" heatid="13018" />
                <RESULT resultid="6142" eventid="15" status="DSQ" swimtime="00:02:49.47" lane="1" heatid="15007" comment="nach der 2. Wende mehrere Delphinkicks.">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:22.43" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1323" birthdate="2014-01-01" gender="F" lastname="Leschinski" firstname="Mariella" license="448018">
              <RESULTS>
                <RESULT resultid="6143" eventid="17" swimtime="00:01:06.69" lane="2" heatid="17005" />
                <RESULT resultid="6144" eventid="19" swimtime="00:00:54.79" lane="3" heatid="19011" />
                <RESULT resultid="6145" eventid="27" swimtime="00:01:06.01" lane="6" heatid="27007" />
                <RESULT resultid="6146" eventid="29" swimtime="00:00:43.57" lane="3" heatid="29009" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1324" birthdate="2014-01-01" gender="F" lastname="Kasielke" firstname="Marlene" license="463191">
              <RESULTS>
                <RESULT resultid="6147" eventid="29" swimtime="00:01:01.23" lane="5" heatid="29001" />
                <RESULT resultid="6148" eventid="31" status="DSQ" swimtime="00:01:31.15" lane="4" heatid="31001" comment="Start vor dem Startsignal." />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1325" birthdate="2014-01-01" gender="F" lastname="Kirsten" firstname="Marta" license="448042">
              <RESULTS>
                <RESULT resultid="6149" eventid="17" swimtime="00:00:55.59" lane="5" heatid="17012" />
                <RESULT resultid="6150" eventid="19" swimtime="00:00:58.05" lane="3" heatid="19006" />
                <RESULT resultid="6151" eventid="25" swimtime="00:00:47.05" lane="8" heatid="25019" />
                <RESULT resultid="6152" eventid="29" swimtime="00:00:43.17" lane="7" heatid="29010" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1326" birthdate="2014-01-01" gender="M" lastname="Warstat" firstname="Mateo" license="463190">
              <RESULTS>
                <RESULT resultid="6153" eventid="18" swimtime="00:01:04.23" lane="3" heatid="18007" />
                <RESULT resultid="6154" eventid="22" swimtime="00:01:05.73" lane="3" heatid="22006" />
                <RESULT resultid="6155" eventid="26" swimtime="00:00:57.56" lane="1" heatid="26003" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1327" birthdate="2008-01-01" gender="F" lastname="Brendler" firstname="Mathilde" license="380792">
              <RESULTS>
                <RESULT resultid="6156" eventid="5" swimtime="00:00:36.40" lane="3" heatid="5008" />
                <RESULT resultid="6157" eventid="10" swimtime="00:01:24.89" lane="6" heatid="10013" />
                <RESULT resultid="6158" eventid="19" swimtime="00:00:46.45" lane="6" heatid="19021" />
                <RESULT resultid="6159" eventid="25" swimtime="00:00:37.94" lane="8" heatid="25032" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1328" birthdate="2007-01-01" gender="F" lastname="Schubert" firstname="Mattea" license="380811">
              <RESULTS>
                <RESULT resultid="6160" eventid="5" swimtime="00:00:28.86" lane="5" heatid="5014" />
                <RESULT resultid="6161" eventid="12" swimtime="00:00:26.61" lane="4" heatid="12018" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1329" birthdate="2015-01-01" gender="M" lastname="Kolkowski" firstname="Max" license="463197">
              <RESULTS>
                <RESULT resultid="6162" eventid="18" status="DSQ" swimtime="00:01:08.60" lane="5" heatid="18005" comment="Start vor dem Startsignal." />
                <RESULT resultid="6163" eventid="20" swimtime="00:01:02.54" lane="5" heatid="20004" />
                <RESULT resultid="6164" eventid="26" swimtime="00:00:56.48" lane="2" heatid="26005" />
                <RESULT resultid="6165" eventid="30" swimtime="00:00:49.56" lane="8" heatid="30004" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1330" birthdate="2011-01-01" gender="M" lastname="Schwarzlose" firstname="Max" license="424896">
              <RESULTS>
                <RESULT resultid="6166" eventid="20" swimtime="00:00:45.50" lane="5" heatid="20014" />
                <RESULT resultid="6167" eventid="26" swimtime="00:00:40.83" lane="1" heatid="26019" />
                <RESULT resultid="6168" eventid="34" swimtime="00:01:24.52" lane="3" heatid="34007" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1331" birthdate="2011-01-01" gender="M" lastname="Bauer" firstname="Maximilian" license="433488">
              <RESULTS>
                <RESULT resultid="6169" eventid="20" status="WDR" swimtime="00:00:00.00" lane="6" heatid="20011" />
                <RESULT resultid="6170" eventid="26" status="WDR" swimtime="00:00:00.00" lane="5" heatid="26008" />
                <RESULT resultid="6171" eventid="34" status="WDR" swimtime="00:00:00.00" lane="8" heatid="34002" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1332" birthdate="2015-01-01" gender="F" lastname="Stange" firstname="Merle" license="463204">
              <RESULTS>
                <RESULT resultid="6172" eventid="17" swimtime="00:01:15.48" lane="4" heatid="17007" />
                <RESULT resultid="6173" eventid="19" swimtime="00:01:09.98" lane="7" heatid="19002" />
                <RESULT resultid="6174" eventid="25" swimtime="00:00:59.29" lane="4" heatid="25007" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1333" birthdate="2012-01-01" gender="F" lastname="Schramm" firstname="Mia" license="436911">
              <RESULTS>
                <RESULT resultid="6175" eventid="3" swimtime="00:01:44.62" lane="5" heatid="3004" />
                <RESULT resultid="6176" eventid="5" swimtime="00:00:45.72" lane="1" heatid="5004" />
                <RESULT resultid="6177" eventid="10" swimtime="00:01:38.91" lane="7" heatid="10006" />
                <RESULT resultid="6178" eventid="14" status="DSQ" swimtime="00:03:38.63" lane="4" heatid="14002" comment="Start vor dem Startsignal.">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:46.71" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="6179" eventid="19" swimtime="00:00:49.03" lane="7" heatid="19017" />
                <RESULT resultid="6180" eventid="27" swimtime="00:01:04.31" lane="6" heatid="27008" />
                <RESULT resultid="6181" eventid="31" swimtime="00:01:00.42" lane="5" heatid="31001" />
                <RESULT resultid="6182" eventid="37" swimtime="00:03:28.16" lane="3" heatid="37002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:43.50" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1334" birthdate="2012-01-01" gender="M" lastname="Martin" firstname="Mika-Frederik" license="436899">
              <RESULTS>
                <RESULT resultid="6183" eventid="6" swimtime="00:00:30.46" lane="2" heatid="6010" />
                <RESULT resultid="6184" eventid="13" swimtime="00:00:29.43" lane="6" heatid="13015" />
                <RESULT resultid="6185" eventid="26" swimtime="00:00:34.07" lane="3" heatid="26023" />
                <RESULT resultid="6186" eventid="36" swimtime="00:01:09.42" lane="7" heatid="36003" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1335" birthdate="2008-01-01" gender="F" lastname="Junge" firstname="Miriam" license="390588">
              <RESULTS>
                <RESULT resultid="6187" eventid="3" swimtime="00:01:36.73" lane="8" heatid="3009" />
                <RESULT resultid="6188" eventid="12" status="DSQ" swimtime="00:00:34.54" lane="5" heatid="12010" comment="Start vor dem Startsignal." />
                <RESULT resultid="6189" eventid="14" swimtime="00:03:25.77" lane="4" heatid="14005">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:40.79" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="6190" eventid="19" swimtime="00:00:44.67" lane="5" heatid="19022" />
                <RESULT resultid="6191" eventid="33" swimtime="00:01:17.80" lane="1" heatid="33012" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1336" birthdate="2014-01-01" gender="F" lastname="Rudolph" firstname="Nienke" license="448172">
              <RESULTS>
                <RESULT resultid="6192" eventid="17" swimtime="00:00:57.84" lane="5" heatid="17009" />
                <RESULT resultid="6193" eventid="19" swimtime="00:00:56.69" lane="4" heatid="19014" />
                <RESULT resultid="6194" eventid="25" swimtime="00:00:47.26" lane="6" heatid="25018" />
                <RESULT resultid="6195" eventid="27" swimtime="00:01:05.93" lane="3" heatid="27006" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1337" birthdate="2013-01-01" gender="M" lastname="Wiese" firstname="Niklas" license="445789">
              <RESULTS>
                <RESULT resultid="6196" eventid="4" swimtime="00:01:45.29" lane="2" heatid="4006" />
                <RESULT resultid="6197" eventid="11" swimtime="00:01:35.51" lane="4" heatid="11006" />
                <RESULT resultid="6198" eventid="13" swimtime="00:00:38.86" lane="1" heatid="13005" />
                <RESULT resultid="6199" eventid="20" swimtime="00:00:48.76" lane="1" heatid="20014" />
                <RESULT resultid="6200" eventid="26" swimtime="00:00:43.11" lane="2" heatid="26017" />
                <RESULT resultid="6201" eventid="28" swimtime="00:01:02.34" lane="8" heatid="28007" />
                <RESULT resultid="6202" eventid="34" swimtime="00:01:26.35" lane="3" heatid="34006" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1338" birthdate="2015-01-01" gender="M" lastname="Suha" firstname="Noah" license="463194">
              <RESULTS>
                <RESULT resultid="6203" eventid="20" swimtime="00:01:03.32" lane="1" heatid="20003" />
                <RESULT resultid="6204" eventid="22" swimtime="00:01:20.51" lane="2" heatid="22002" />
                <RESULT resultid="6205" eventid="26" swimtime="00:00:57.27" lane="1" heatid="26005" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1339" birthdate="2015-01-01" gender="M" lastname="Mattke" firstname="Pepe Luis" license="463212">
              <RESULTS>
                <RESULT resultid="6206" eventid="18" swimtime="00:01:17.78" lane="5" heatid="18004" />
                <RESULT resultid="6207" eventid="22" swimtime="00:01:10.63" lane="4" heatid="22003" />
                <RESULT resultid="6208" eventid="26" swimtime="00:00:54.87" lane="8" heatid="26007" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1340" birthdate="2011-01-01" gender="M" lastname="Schulze" firstname="Philipp" license="433489">
              <RESULTS>
                <RESULT resultid="6209" eventid="4" swimtime="00:02:07.60" lane="8" heatid="4002" />
                <RESULT resultid="6210" eventid="13" swimtime="00:00:45.25" lane="7" heatid="13002" />
                <RESULT resultid="6211" eventid="15" swimtime="00:04:37.60" lane="1" heatid="15002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:02:17.28" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1341" birthdate="2014-01-01" gender="F" lastname="Müller" firstname="Pia" license="448027">
              <RESULTS>
                <RESULT resultid="6212" eventid="17" swimtime="00:01:08.29" lane="6" heatid="17004" />
                <RESULT resultid="6213" eventid="21" swimtime="00:01:00.65" lane="1" heatid="21005" />
                <RESULT resultid="6214" eventid="25" swimtime="00:00:48.32" lane="5" heatid="25013" />
                <RESULT resultid="6215" eventid="29" swimtime="00:00:41.35" lane="8" heatid="29012" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1342" birthdate="2014-01-01" gender="M" lastname="Glaser" firstname="Raphael" license="448022">
              <RESULTS>
                <RESULT resultid="6216" eventid="18" swimtime="00:00:58.95" lane="5" heatid="18009" />
                <RESULT resultid="6217" eventid="20" swimtime="00:00:57.13" lane="2" heatid="20006" />
                <RESULT resultid="6218" eventid="26" swimtime="00:00:49.61" lane="3" heatid="26008" />
                <RESULT resultid="6219" eventid="30" swimtime="00:00:43.68" lane="1" heatid="30005" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1343" birthdate="2010-01-01" gender="M" lastname="Zesewitz" firstname="Raphael" license="412733">
              <RESULTS>
                <RESULT resultid="6220" eventid="2" swimtime="00:02:31.01" lane="6" heatid="2008">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:12.95" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="6221" eventid="9" swimtime="00:02:40.62" lane="5" heatid="9001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:14.98" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1344" birthdate="2012-01-01" gender="M" lastname="Petzold" firstname="Richard" license="445370">
              <RESULTS>
                <RESULT resultid="6222" eventid="20" status="WDR" swimtime="00:00:00.00" lane="2" heatid="20009" />
                <RESULT resultid="6223" eventid="26" status="WDR" swimtime="00:00:00.00" lane="8" heatid="26012" />
                <RESULT resultid="6224" eventid="28" status="WDR" swimtime="00:00:00.00" lane="2" heatid="28003" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1345" birthdate="2015-01-01" gender="M" lastname="Franke" firstname="Robin" license="463214">
              <RESULTS>
                <RESULT resultid="6225" eventid="20" swimtime="00:01:04.23" lane="8" heatid="20003" />
                <RESULT resultid="6226" eventid="22" swimtime="00:01:17.48" lane="3" heatid="22002" />
                <RESULT resultid="6227" eventid="26" swimtime="00:01:02.90" lane="2" heatid="26003" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1346" birthdate="2015-01-01" gender="F" lastname="Fritzsche" firstname="Sara" license="463219">
              <RESULTS>
                <RESULT resultid="6228" eventid="17" swimtime="00:01:10.84" lane="3" heatid="17006" />
                <RESULT resultid="6229" eventid="19" swimtime="00:01:10.38" lane="3" heatid="19003" />
                <RESULT resultid="6230" eventid="25" swimtime="00:01:01.44" lane="5" heatid="25004" />
                <RESULT resultid="6231" eventid="27" swimtime="00:01:15.82" lane="4" heatid="27003" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1347" birthdate="2012-01-01" gender="F" lastname="Schellhammer" firstname="Sarafina" license="444321">
              <RESULTS>
                <RESULT resultid="6232" eventid="3" swimtime="00:01:37.83" lane="4" heatid="3008" />
                <RESULT resultid="6233" eventid="5" swimtime="00:00:41.29" lane="7" heatid="5006" />
                <RESULT resultid="6234" eventid="23" swimtime="00:02:57.89" lane="5" heatid="23005">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:25.34" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="6235" eventid="27" swimtime="00:00:56.33" lane="7" heatid="27011" />
                <RESULT resultid="6236" eventid="33" swimtime="00:01:22.17" lane="6" heatid="33013" />
                <RESULT resultid="6237" eventid="37" swimtime="00:03:04.42" lane="2" heatid="37006">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:31.49" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1348" birthdate="2014-01-01" gender="M" lastname="Körner" firstname="Simon Friedrich" license="464255">
              <RESULTS>
                <RESULT resultid="6238" eventid="18" swimtime="00:01:05.74" lane="6" heatid="18008" />
                <RESULT resultid="6239" eventid="20" swimtime="00:00:59.08" lane="7" heatid="20004" />
                <RESULT resultid="6240" eventid="22" swimtime="00:00:59.65" lane="7" heatid="22007" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1349" birthdate="2014-01-01" gender="M" lastname="Sperling" firstname="Sirko" license="452436">
              <RESULTS>
                <RESULT resultid="6241" eventid="18" swimtime="00:01:01.84" lane="1" heatid="18005" />
                <RESULT resultid="6242" eventid="22" swimtime="00:00:57.29" lane="2" heatid="22008" />
                <RESULT resultid="6243" eventid="28" swimtime="00:01:04.95" lane="1" heatid="28004" />
                <RESULT resultid="6244" eventid="30" swimtime="00:00:36.39" lane="5" heatid="30008" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1350" birthdate="2011-01-01" gender="F" lastname="Abdel Bary" firstname="Soraya" license="424559">
              <RESULTS>
                <RESULT resultid="6245" eventid="3" status="WDR" swimtime="00:00:00.00" lane="7" heatid="3003" />
                <RESULT resultid="6246" eventid="5" status="WDR" swimtime="00:00:00.00" lane="4" heatid="5002" />
                <RESULT resultid="6247" eventid="12" status="WDR" swimtime="00:00:00.00" lane="6" heatid="12005" />
                <RESULT resultid="6248" eventid="14" status="WDR" swimtime="00:00:00.00" lane="2" heatid="14003" />
                <RESULT resultid="6249" eventid="19" status="WDR" swimtime="00:00:00.00" lane="6" heatid="19019" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1351" birthdate="2015-01-01" gender="M" lastname="Schweigler" firstname="Theo" license="463203">
              <RESULTS>
                <RESULT resultid="6250" eventid="20" status="WDR" swimtime="00:00:00.00" lane="5" heatid="20001" />
                <RESULT resultid="6251" eventid="26" status="WDR" swimtime="00:00:00.00" lane="3" heatid="26004" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1352" birthdate="2012-01-01" gender="M" lastname="Neumann" firstname="Till" license="436908">
              <RESULTS>
                <RESULT resultid="6252" eventid="20" swimtime="00:00:50.26" lane="5" heatid="20010" />
                <RESULT resultid="6253" eventid="26" swimtime="00:00:49.14" lane="4" heatid="26013" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1353" birthdate="2014-01-01" gender="M" lastname="Müller" firstname="Tristan" license="448066">
              <RESULTS>
                <RESULT resultid="6254" eventid="18" swimtime="00:01:18.20" lane="8" heatid="18003" />
                <RESULT resultid="6255" eventid="20" swimtime="00:00:56.24" lane="3" heatid="20005" />
                <RESULT resultid="6256" eventid="26" swimtime="00:00:59.30" lane="4" heatid="26003" />
                <RESULT resultid="6257" eventid="30" swimtime="00:00:46.65" lane="4" heatid="30003" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1354" birthdate="2013-01-01" gender="M" lastname="Paris" firstname="Yanic" license="448044">
              <RESULTS>
                <RESULT resultid="6258" eventid="2" swimtime="00:03:31.92" lane="5" heatid="2003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:37.69" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="6259" eventid="6" swimtime="00:00:42.44" lane="2" heatid="6004" />
                <RESULT resultid="6260" eventid="11" swimtime="00:01:34.51" lane="8" heatid="11006" />
                <RESULT resultid="6261" eventid="13" swimtime="00:00:38.68" lane="4" heatid="13003" />
                <RESULT resultid="6262" eventid="20" swimtime="00:00:50.22" lane="7" heatid="20012" />
                <RESULT resultid="6263" eventid="26" swimtime="00:00:43.10" lane="5" heatid="26015" />
                <RESULT resultid="6264" eventid="32" swimtime="00:00:59.19" lane="6" heatid="32002" />
                <RESULT resultid="6265" eventid="38" swimtime="00:03:19.58" lane="5" heatid="38001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:38.99" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY number="1" gender="X" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="5821" eventid="7" swimtime="00:02:09.45" lane="4" heatid="7003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:09.63" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1343" number="1" />
                    <RELAYPOSITION athleteid="1267" number="2" />
                    <RELAYPOSITION athleteid="1320" number="3" />
                    <RELAYPOSITION athleteid="1334" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" gender="X" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="5822" eventid="16" swimtime="00:01:58.07" lane="4" heatid="16002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:03.42" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1322" number="1" />
                    <RELAYPOSITION athleteid="1247" number="2" />
                    <RELAYPOSITION athleteid="1289" number="3" />
                    <RELAYPOSITION athleteid="1328" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="2" gender="X" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="5823" eventid="7" swimtime="00:02:31.62" lane="8" heatid="7003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:21.34" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1314" number="1" />
                    <RELAYPOSITION athleteid="1347" number="2" />
                    <RELAYPOSITION athleteid="1270" number="3" />
                    <RELAYPOSITION athleteid="1298" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="3" gender="X" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="5824" eventid="7" swimtime="00:02:36.47" lane="2" heatid="7002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:23.90" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1292" number="1" />
                    <RELAYPOSITION athleteid="1337" number="2" />
                    <RELAYPOSITION athleteid="1249" number="3" />
                    <RELAYPOSITION athleteid="1272" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="4" gender="X" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="5825" eventid="7" swimtime="00:02:48.94" lane="5" heatid="7001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:31.93" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1259" number="1" />
                    <RELAYPOSITION athleteid="1290" number="2" />
                    <RELAYPOSITION athleteid="1354" number="3" />
                    <RELAYPOSITION athleteid="1269" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="5" gender="X" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="5826" eventid="7" swimtime="00:02:49.43" lane="3" heatid="7001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:33.57" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1303" number="1" />
                    <RELAYPOSITION athleteid="1285" number="2" />
                    <RELAYPOSITION athleteid="1258" number="3" />
                    <RELAYPOSITION athleteid="1260" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB name="FC Erzgebirge Aue" nation="GER" region="12" code="7123">
          <ATHLETES>
            <ATHLETE athleteid="1035" birthdate="2009-01-01" gender="M" lastname="Weber" firstname="Anton" license="395001">
              <RESULTS>
                <RESULT resultid="4804" eventid="4" swimtime="00:01:39.90" lane="7" heatid="4006" />
                <RESULT resultid="4805" eventid="13" swimtime="00:00:32.38" lane="4" heatid="13011" />
                <RESULT resultid="4806" eventid="15" swimtime="00:03:42.70" lane="6" heatid="15003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:49.34" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="4807" eventid="20" swimtime="00:00:45.99" lane="3" heatid="20014" />
                <RESULT resultid="4808" eventid="26" swimtime="00:00:41.57" lane="1" heatid="26014" />
                <RESULT resultid="4809" eventid="34" swimtime="00:01:15.99" lane="8" heatid="34004" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1036" birthdate="2012-01-01" gender="F" lastname="Tenelsen" firstname="Fenja" license="434707">
              <RESULTS>
                <RESULT resultid="4810" eventid="3" swimtime="00:01:42.85" lane="5" heatid="3006" />
                <RESULT resultid="4811" eventid="10" swimtime="00:01:34.69" lane="5" heatid="10009" />
                <RESULT resultid="4812" eventid="12" swimtime="00:00:36.22" lane="6" heatid="12009" />
                <RESULT resultid="4813" eventid="17" swimtime="00:00:55.82" lane="2" heatid="17013" />
                <RESULT resultid="4814" eventid="19" swimtime="00:00:46.81" lane="2" heatid="19019" />
                <RESULT resultid="4815" eventid="25" swimtime="00:00:42.72" lane="5" heatid="25026" />
                <RESULT resultid="4816" eventid="27" swimtime="00:00:57.49" lane="5" heatid="27008" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1037" birthdate="2009-01-01" gender="M" lastname="Grunert" firstname="Ferdinand" license="395006">
              <RESULTS>
                <RESULT resultid="4817" eventid="4" swimtime="00:01:37.32" lane="4" heatid="4006" />
                <RESULT resultid="4818" eventid="6" swimtime="00:00:39.16" lane="7" heatid="6005" />
                <RESULT resultid="4819" eventid="11" swimtime="00:01:34.58" lane="3" heatid="11007" />
                <RESULT resultid="4820" eventid="13" swimtime="00:00:33.59" lane="1" heatid="13010" />
                <RESULT resultid="4821" eventid="20" swimtime="00:00:44.20" lane="1" heatid="20017" />
                <RESULT resultid="4822" eventid="26" swimtime="00:00:43.38" lane="8" heatid="26014" />
                <RESULT resultid="4823" eventid="34" swimtime="00:01:16.51" lane="1" heatid="34010" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1038" birthdate="2012-01-01" gender="M" lastname="Kraus" firstname="Finn" license="432063">
              <RESULTS>
                <RESULT resultid="4824" eventid="4" swimtime="00:01:46.36" lane="3" heatid="4004" />
                <RESULT resultid="4825" eventid="6" swimtime="00:00:48.45" lane="3" heatid="6002" />
                <RESULT resultid="4826" eventid="13" swimtime="00:00:35.66" lane="1" heatid="13008" />
                <RESULT resultid="4827" eventid="20" swimtime="00:00:46.97" lane="5" heatid="20013" />
                <RESULT resultid="4828" eventid="26" swimtime="00:00:40.75" lane="5" heatid="26019" />
                <RESULT resultid="4829" eventid="28" swimtime="00:01:02.90" lane="1" heatid="28007" />
                <RESULT resultid="4830" eventid="34" swimtime="00:01:23.15" lane="7" heatid="34006" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1039" birthdate="2006-01-01" gender="M" lastname="Heydel" firstname="Ian" license="433479">
              <RESULTS>
                <RESULT resultid="4831" eventid="4" swimtime="00:01:25.46" lane="7" heatid="4010" />
                <RESULT resultid="4832" eventid="6" swimtime="00:00:32.97" lane="3" heatid="6009" />
                <RESULT resultid="4833" eventid="13" swimtime="00:00:30.06" lane="5" heatid="13015" />
                <RESULT resultid="4834" eventid="20" swimtime="00:00:38.45" lane="6" heatid="20021" />
                <RESULT resultid="4835" eventid="26" swimtime="00:00:34.45" lane="4" heatid="26023" />
                <RESULT resultid="4836" eventid="34" swimtime="00:01:07.74" lane="2" heatid="34013" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1040" birthdate="2006-01-01" gender="F" lastname="Fritzsch" firstname="Julie" license="363418">
              <RESULTS>
                <RESULT resultid="4837" eventid="3" swimtime="00:01:38.89" lane="3" heatid="3008" />
                <RESULT resultid="4838" eventid="5" swimtime="00:00:39.38" lane="2" heatid="5005" />
                <RESULT resultid="4839" eventid="12" swimtime="00:00:33.44" lane="2" heatid="12014" />
                <RESULT resultid="4840" eventid="19" swimtime="00:00:45.36" lane="2" heatid="19023" />
                <RESULT resultid="4841" eventid="23" swimtime="00:02:43.91" lane="1" heatid="23010">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:16.43" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="4842" eventid="33" swimtime="00:01:13.14" lane="5" heatid="33014" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1041" birthdate="2010-01-01" gender="F" lastname="Sandow" firstname="Kena" license="433481">
              <RESULTS>
                <RESULT resultid="4843" eventid="5" status="DNS" swimtime="00:00:00.00" lane="5" heatid="5007" />
                <RESULT resultid="4844" eventid="10" status="DNS" swimtime="00:00:00.00" lane="3" heatid="10009" />
                <RESULT resultid="4845" eventid="12" status="DNS" swimtime="00:00:00.00" lane="1" heatid="12011" />
                <RESULT resultid="4846" eventid="19" swimtime="00:00:46.11" lane="1" heatid="19019" />
                <RESULT resultid="4847" eventid="25" swimtime="00:00:40.72" lane="1" heatid="25027" />
                <RESULT resultid="4848" eventid="33" swimtime="00:01:18.85" lane="8" heatid="33012" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1042" birthdate="2008-01-01" gender="M" lastname="Ullmann" firstname="Konstantin" license="349898">
              <RESULTS>
                <RESULT resultid="4849" eventid="4" swimtime="00:01:27.63" lane="1" heatid="4004" />
                <RESULT resultid="4850" eventid="6" swimtime="00:00:30.75" lane="5" heatid="6010" />
                <RESULT resultid="4851" eventid="11" swimtime="00:01:16.70" lane="8" heatid="11012" />
                <RESULT resultid="4852" eventid="13" swimtime="00:00:28.96" lane="6" heatid="13017" />
                <RESULT resultid="4853" eventid="20" swimtime="00:00:38.39" lane="5" heatid="20020" />
                <RESULT resultid="4854" eventid="26" swimtime="00:00:32.71" lane="7" heatid="26024" />
                <RESULT resultid="4855" eventid="34" swimtime="00:01:03.92" lane="7" heatid="34014" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1043" birthdate="2012-01-01" gender="F" lastname="Riediger" firstname="Lani" license="459623">
              <RESULTS>
                <RESULT resultid="4856" eventid="3" status="DSQ" swimtime="00:01:45.66" lane="1" heatid="3006" comment="Beine auf der zweiten Bahn nicht gleichzeitig bewegt." />
                <RESULT resultid="4857" eventid="5" swimtime="00:00:52.24" lane="3" heatid="5002" />
                <RESULT resultid="4858" eventid="12" swimtime="00:00:37.63" lane="2" heatid="12007" />
                <RESULT resultid="4859" eventid="19" swimtime="00:00:47.21" lane="4" heatid="19019" />
                <RESULT resultid="4860" eventid="25" status="DSQ" swimtime="00:00:43.13" lane="3" heatid="25020" comment="Start vor dem Startsignal." />
                <RESULT resultid="4861" eventid="27" status="DSQ" swimtime="00:00:57.17" lane="3" heatid="27012" comment="Beine nicht gleichzeitig bewegt." />
                <RESULT resultid="4862" eventid="33" swimtime="00:01:24.67" lane="5" heatid="33007" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1044" birthdate="2011-01-01" gender="F" lastname="Weidauer" firstname="Lavinia" license="419465">
              <RESULTS>
                <RESULT resultid="4863" eventid="3" swimtime="00:01:43.39" lane="8" heatid="3005" />
                <RESULT resultid="4864" eventid="5" swimtime="00:00:37.96" lane="4" heatid="5007" />
                <RESULT resultid="4865" eventid="10" swimtime="00:01:30.56" lane="1" heatid="10010" />
                <RESULT resultid="4866" eventid="12" swimtime="00:00:33.04" lane="5" heatid="12012" />
                <RESULT resultid="4867" eventid="19" swimtime="00:00:45.77" lane="7" heatid="19019" />
                <RESULT resultid="4868" eventid="25" swimtime="00:00:39.59" lane="5" heatid="25030" />
                <RESULT resultid="4869" eventid="33" swimtime="00:01:14.55" lane="4" heatid="33011" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1045" birthdate="2012-01-01" gender="F" lastname="Nitsche" firstname="Lea" license="459626">
              <RESULTS>
                <RESULT resultid="4870" eventid="3" swimtime="00:01:51.72" lane="8" heatid="3004" />
                <RESULT resultid="4871" eventid="5" swimtime="00:00:50.52" lane="5" heatid="5002" />
                <RESULT resultid="4872" eventid="10" swimtime="00:01:44.02" lane="1" heatid="10003" />
                <RESULT resultid="4873" eventid="12" swimtime="00:00:39.81" lane="4" heatid="12006" />
                <RESULT resultid="4874" eventid="19" swimtime="00:00:50.50" lane="5" heatid="19014" />
                <RESULT resultid="4875" eventid="27" swimtime="00:00:59.39" lane="2" heatid="27012" />
                <RESULT resultid="4876" eventid="33" swimtime="00:01:35.01" lane="7" heatid="33005" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1046" birthdate="2010-01-01" gender="F" lastname="Ullmann" firstname="Linn" license="419258">
              <RESULTS>
                <RESULT resultid="4877" eventid="3" swimtime="00:01:33.30" lane="6" heatid="3009" />
                <RESULT resultid="4878" eventid="10" swimtime="00:01:37.54" lane="4" heatid="10006" />
                <RESULT resultid="4879" eventid="12" swimtime="00:00:35.30" lane="6" heatid="12010" />
                <RESULT resultid="4880" eventid="14" swimtime="00:03:25.31" lane="6" heatid="14006">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:38.83" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="4881" eventid="19" swimtime="00:00:43.35" lane="3" heatid="19024" />
                <RESULT resultid="4882" eventid="25" swimtime="00:00:42.16" lane="7" heatid="25026" />
                <RESULT resultid="4883" eventid="33" swimtime="00:01:18.99" lane="3" heatid="33010" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1047" birthdate="2009-01-01" gender="F" lastname="Petrick" firstname="Martha" license="433480">
              <RESULTS>
                <RESULT resultid="4884" eventid="3" swimtime="00:01:32.69" lane="7" heatid="3009" />
                <RESULT resultid="4885" eventid="5" swimtime="00:00:37.09" lane="5" heatid="5009" />
                <RESULT resultid="4886" eventid="12" swimtime="00:00:32.76" lane="3" heatid="12015" />
                <RESULT resultid="4887" eventid="19" swimtime="00:00:42.67" lane="2" heatid="19024" />
                <RESULT resultid="4888" eventid="25" swimtime="00:00:38.43" lane="6" heatid="25032" />
                <RESULT resultid="4889" eventid="33" swimtime="00:01:10.85" lane="8" heatid="33017" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1048" birthdate="2010-01-01" gender="M" lastname="Wietz" firstname="Paul" license="395002">
              <RESULTS>
                <RESULT resultid="4890" eventid="4" swimtime="00:01:43.53" lane="6" heatid="4004" />
                <RESULT resultid="4891" eventid="6" swimtime="00:00:48.56" lane="3" heatid="6003" />
                <RESULT resultid="4892" eventid="13" swimtime="00:00:34.98" lane="1" heatid="13011" />
                <RESULT resultid="4893" eventid="20" swimtime="00:00:47.05" lane="8" heatid="20015" />
                <RESULT resultid="4894" eventid="24" swimtime="00:02:50.04" lane="2" heatid="24006">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:19.55" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="4895" eventid="26" swimtime="00:00:41.50" lane="1" heatid="26021" />
                <RESULT resultid="4896" eventid="34" swimtime="00:01:15.67" lane="5" heatid="34010" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1049" birthdate="2011-01-01" gender="M" lastname="Lötzsch" firstname="Theo" license="419466">
              <RESULTS>
                <RESULT resultid="4897" eventid="4" swimtime="00:01:50.85" lane="2" heatid="4004" />
                <RESULT resultid="4898" eventid="11" swimtime="00:01:39.37" lane="6" heatid="11005" />
                <RESULT resultid="4899" eventid="13" swimtime="00:00:36.99" lane="3" heatid="13007" />
                <RESULT resultid="4900" eventid="15" swimtime="00:03:59.86" lane="8" heatid="15003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:57.46" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="4901" eventid="20" swimtime="00:00:49.90" lane="4" heatid="20011" />
                <RESULT resultid="4902" eventid="26" swimtime="00:00:44.32" lane="4" heatid="26014" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1050" birthdate="2008-01-01" gender="M" lastname="Kraus" firstname="Tim" license="395174">
              <RESULTS>
                <RESULT resultid="4903" eventid="4" swimtime="00:01:33.64" lane="5" heatid="4008" />
                <RESULT resultid="4904" eventid="6" swimtime="00:00:37.39" lane="6" heatid="6002" />
                <RESULT resultid="4905" eventid="11" swimtime="00:01:21.61" lane="5" heatid="11009" />
                <RESULT resultid="4906" eventid="13" swimtime="00:00:28.51" lane="4" heatid="13016" />
                <RESULT resultid="4907" eventid="20" swimtime="00:00:41.99" lane="1" heatid="20019" />
                <RESULT resultid="4908" eventid="26" swimtime="00:00:34.97" lane="8" heatid="26023" />
                <RESULT resultid="4909" eventid="34" swimtime="00:01:07.19" lane="1" heatid="34013" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1051" birthdate="2012-01-01" gender="F" lastname="Müller" firstname="Zoe" license="417100">
              <RESULTS>
                <RESULT resultid="4910" eventid="5" swimtime="00:00:45.91" lane="8" heatid="5004" />
                <RESULT resultid="4911" eventid="10" swimtime="00:01:27.63" lane="4" heatid="10012" />
                <RESULT resultid="4912" eventid="12" swimtime="00:00:36.21" lane="3" heatid="12009" />
                <RESULT resultid="4913" eventid="21" swimtime="00:00:54.81" lane="2" heatid="21013" />
                <RESULT resultid="4914" eventid="25" swimtime="00:00:39.86" lane="7" heatid="25030" />
                <RESULT resultid="4915" eventid="31" swimtime="00:00:55.93" lane="7" heatid="31004" />
                <RESULT resultid="4916" eventid="37" swimtime="00:03:05.81" lane="7" heatid="37006">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:30.54" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY number="1" gender="X" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="4801" eventid="16" swimtime="00:02:16.43" lane="7" heatid="16002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:16.39" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1047" number="1" />
                    <RELAYPOSITION athleteid="1039" number="2" />
                    <RELAYPOSITION athleteid="1042" number="3" />
                    <RELAYPOSITION athleteid="1050" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" gender="X" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="4802" eventid="7" swimtime="00:02:42.93" lane="7" heatid="7002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:24.58" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1051" number="1" />
                    <RELAYPOSITION athleteid="1046" number="2" />
                    <RELAYPOSITION athleteid="1048" number="3" />
                    <RELAYPOSITION athleteid="1044" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="2" gender="X" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="4803" eventid="7" swimtime="00:02:56.99" lane="8" heatid="7002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:32.64" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1049" number="1" />
                    <RELAYPOSITION athleteid="1036" number="2" />
                    <RELAYPOSITION athleteid="1038" number="3" />
                    <RELAYPOSITION athleteid="1043" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB name="Post SV Dresden" nation="GER" region="12" code="3348">
          <ATHLETES>
            <ATHLETE athleteid="1061" birthdate="2006-01-01" gender="F" lastname="Siemens" firstname="Alice" license="402495">
              <RESULTS>
                <RESULT resultid="4960" eventid="19" swimtime="00:00:48.08" lane="6" heatid="19020" />
                <RESULT resultid="4961" eventid="23" swimtime="00:02:51.92" lane="4" heatid="23004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:21.58" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="4962" eventid="33" swimtime="00:01:16.94" lane="3" heatid="33013" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1062" birthdate="2009-01-01" gender="F" lastname="Belling" firstname="Caroline" license="417614">
              <RESULTS>
                <RESULT resultid="4963" eventid="23" swimtime="00:02:50.28" lane="8" heatid="23006">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:23.28" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="4964" eventid="25" swimtime="00:00:38.91" lane="2" heatid="25024" />
                <RESULT resultid="4965" eventid="33" swimtime="00:01:16.51" lane="7" heatid="33012" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1063" birthdate="2006-01-01" gender="F" lastname="Specht" firstname="Franziska" license="349837">
              <RESULTS>
                <RESULT resultid="4966" eventid="23" swimtime="00:02:27.19" lane="6" heatid="23009">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:08.06" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="4967" eventid="25" swimtime="00:00:33.84" lane="5" heatid="25034" />
                <RESULT resultid="4968" eventid="33" swimtime="00:01:06.42" lane="8" heatid="33018" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1064" birthdate="2010-01-01" gender="F" lastname="Leibling" firstname="Janka" license="431463">
              <RESULTS>
                <RESULT resultid="4969" eventid="19" status="DSQ" swimtime="00:00:44.66" lane="3" heatid="19022" comment="Start vor dem Startsignal." />
                <RESULT resultid="4970" eventid="23" swimtime="00:02:55.90" lane="3" heatid="23003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:26.14" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="4971" eventid="25" swimtime="00:00:40.34" lane="3" heatid="25025" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1065" birthdate="2007-01-01" gender="F" lastname="Schulze" firstname="Lilly Vivien" license="374475">
              <RESULTS>
                <RESULT resultid="4972" eventid="19" status="WDR" swimtime="00:00:00.00" lane="4" heatid="19022" />
                <RESULT resultid="4973" eventid="23" status="WDR" swimtime="00:00:00.00" lane="5" heatid="23003" />
                <RESULT resultid="4974" eventid="25" status="WDR" swimtime="00:00:00.00" lane="3" heatid="25028" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1066" birthdate="2006-01-01" gender="F" lastname="Würschig" firstname="Mareike" license="335967">
              <RESULTS>
                <RESULT resultid="4975" eventid="23" swimtime="00:03:10.95" lane="1" heatid="23002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:31.56" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="4976" eventid="25" swimtime="00:00:42.47" lane="3" heatid="25026" />
                <RESULT resultid="4977" eventid="33" swimtime="00:01:22.91" lane="3" heatid="33009" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1067" birthdate="2009-01-01" gender="F" lastname="Schukoff" firstname="Melina" license="417613">
              <RESULTS>
                <RESULT resultid="4978" eventid="19" swimtime="00:00:43.42" lane="2" heatid="19026" />
                <RESULT resultid="4979" eventid="23" swimtime="00:02:53.15" lane="1" heatid="23005">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:24.00" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="4980" eventid="25" swimtime="00:00:39.48" lane="7" heatid="25027" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="Post SV Leipzig e.V." nation="GER" region="12" code="3351">
          <ATHLETES>
            <ATHLETE athleteid="332" birthdate="2012-01-01" gender="F" lastname="Schulze" firstname="Zazou" license="440958">
              <RESULTS>
                <RESULT resultid="1600" eventid="3" swimtime="00:01:40.65" lane="5" heatid="3005" />
                <RESULT resultid="1599" eventid="10" status="DSQ" swimtime="00:01:36.02" lane="4" heatid="10008" comment="Start vor dem Startsignal." />
                <RESULT resultid="1598" eventid="12" swimtime="00:00:36.10" lane="2" heatid="12008" />
                <RESULT resultid="1597" eventid="17" swimtime="00:00:53.27" lane="8" heatid="17015" />
                <RESULT resultid="1596" eventid="25" swimtime="00:00:40.51" lane="3" heatid="25027" />
                <RESULT resultid="1595" eventid="37" swimtime="00:03:15.17" lane="1" heatid="37003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:36.17" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="333" birthdate="2014-01-01" gender="M" lastname="Severyuk" firstname="Vincent" license="448125">
              <RESULTS>
                <RESULT resultid="1605" eventid="18" swimtime="00:01:05.98" lane="5" heatid="18008" />
                <RESULT resultid="1604" eventid="22" swimtime="00:01:00.14" lane="4" heatid="22009" />
                <RESULT resultid="1603" eventid="26" swimtime="00:00:50.04" lane="2" heatid="26013" />
                <RESULT resultid="1602" eventid="30" swimtime="00:00:42.39" lane="2" heatid="30008" />
                <RESULT resultid="1601" eventid="34" swimtime="00:01:41.46" lane="8" heatid="34003" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="334" birthdate="2012-01-01" gender="F" lastname="Schindler" firstname="Rosa" license="440950">
              <RESULTS>
                <RESULT resultid="1611" eventid="5" swimtime="00:00:39.66" lane="3" heatid="5007" />
                <RESULT resultid="1610" eventid="10" swimtime="00:01:30.83" lane="7" heatid="10011" />
                <RESULT resultid="1609" eventid="12" swimtime="00:00:36.16" lane="4" heatid="12010" />
                <RESULT resultid="1608" eventid="21" swimtime="00:00:53.90" lane="3" heatid="21013" />
                <RESULT resultid="1607" eventid="25" swimtime="00:00:40.73" lane="7" heatid="25032" />
                <RESULT resultid="1606" eventid="37" status="DSQ" swimtime="00:03:06.96" lane="1" heatid="37006" comment="Bei der 2. Wende wurde die Wende nicht unverzüglich nach Einnahme der Bauchlage ausgeführt.">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:33.80" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="335" birthdate="2012-01-01" gender="F" lastname="Hacker" firstname="Mara" license="440971">
              <RESULTS>
                <RESULT resultid="1617" eventid="5" swimtime="00:00:39.23" lane="6" heatid="5006" />
                <RESULT resultid="1616" eventid="10" swimtime="00:01:32.17" lane="2" heatid="10007" />
                <RESULT resultid="1615" eventid="12" swimtime="00:00:35.36" lane="6" heatid="12008" />
                <RESULT resultid="1614" eventid="17" swimtime="00:01:00.93" lane="5" heatid="17013" />
                <RESULT resultid="1613" eventid="23" swimtime="00:02:59.76" lane="5" heatid="23004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:25.31" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1612" eventid="33" swimtime="00:01:19.41" lane="7" heatid="33010" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="336" birthdate="2014-01-01" gender="M" lastname="Twal" firstname="Malik" license="461707">
              <RESULTS>
                <RESULT resultid="1621" eventid="20" swimtime="00:00:51.44" lane="2" heatid="20011" />
                <RESULT resultid="1620" eventid="28" swimtime="00:01:07.09" lane="6" heatid="28004" />
                <RESULT resultid="1619" eventid="30" swimtime="00:00:45.71" lane="3" heatid="30007" />
                <RESULT resultid="1618" eventid="34" swimtime="00:01:42.08" lane="1" heatid="34003" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="337" birthdate="2013-01-01" gender="M" lastname="Schlegel" firstname="Levi Anton" license="444301">
              <RESULTS>
                <RESULT resultid="1627" eventid="4" swimtime="00:01:48.95" lane="2" heatid="4005" />
                <RESULT resultid="1626" eventid="11" swimtime="00:01:42.12" lane="5" heatid="11002" />
                <RESULT resultid="1625" eventid="15" swimtime="00:03:52.66" lane="6" heatid="15002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:55.61" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1624" eventid="20" swimtime="00:00:50.80" lane="8" heatid="20012" />
                <RESULT resultid="1623" eventid="22" swimtime="00:00:53.73" lane="2" heatid="22009" />
                <RESULT resultid="1622" eventid="28" swimtime="00:00:56.00" lane="4" heatid="28007" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="338" birthdate="2013-01-01" gender="M" lastname="Richter" firstname="Justus" license="444299">
              <RESULTS>
                <RESULT resultid="1633" eventid="4" swimtime="00:01:39.97" lane="4" heatid="4007" />
                <RESULT resultid="1632" eventid="13" swimtime="00:00:38.62" lane="2" heatid="13005" />
                <RESULT resultid="1631" eventid="15" swimtime="00:03:29.59" lane="6" heatid="15004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:43.14" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1630" eventid="20" swimtime="00:00:45.25" lane="8" heatid="20017" />
                <RESULT resultid="1629" eventid="28" swimtime="00:00:55.57" lane="1" heatid="28008" />
                <RESULT resultid="1628" eventid="38" swimtime="00:03:15.65" lane="7" heatid="38003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:36.57" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="339" birthdate="2014-01-01" gender="F" lastname="Hoppe" firstname="Hannah" license="448122">
              <RESULTS>
                <RESULT resultid="1638" eventid="17" swimtime="00:00:59.26" lane="6" heatid="17011" />
                <RESULT resultid="1637" eventid="19" swimtime="00:00:53.06" lane="3" heatid="19015" />
                <RESULT resultid="1636" eventid="25" swimtime="00:00:48.64" lane="1" heatid="25019" />
                <RESULT resultid="1635" eventid="29" swimtime="00:00:41.98" lane="7" heatid="29012" />
                <RESULT resultid="1634" eventid="31" swimtime="00:01:01.28" lane="1" heatid="31005" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="340" birthdate="2014-01-01" gender="F" lastname="Meißner" firstname="Frida" license="448123">
              <RESULTS>
                <RESULT resultid="1643" eventid="17" swimtime="00:00:48.42" lane="5" heatid="17016" />
                <RESULT resultid="1642" eventid="21" swimtime="00:00:48.81" lane="4" heatid="21014" />
                <RESULT resultid="1641" eventid="25" swimtime="00:00:43.32" lane="6" heatid="25025" />
                <RESULT resultid="1640" eventid="29" swimtime="00:00:37.20" lane="5" heatid="29013" />
                <RESULT resultid="1639" eventid="31" swimtime="00:00:53.46" lane="6" heatid="31007" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="341" birthdate="2012-01-01" gender="F" lastname="Waizmann" firstname="Emilia" license="442586">
              <RESULTS>
                <RESULT resultid="1648" eventid="3" swimtime="00:01:53.36" lane="2" heatid="3003" />
                <RESULT resultid="1647" eventid="12" swimtime="00:00:41.93" lane="4" heatid="12003" />
                <RESULT resultid="1646" eventid="21" swimtime="00:00:56.64" lane="1" heatid="21013" />
                <RESULT resultid="1645" eventid="27" swimtime="00:01:02.79" lane="3" heatid="27008" />
                <RESULT resultid="1644" eventid="31" swimtime="00:01:07.56" lane="4" heatid="31002" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="342" birthdate="2012-01-01" gender="F" lastname="Scheel" firstname="Charlotte Luise" license="443056">
              <RESULTS>
                <RESULT resultid="1654" eventid="5" swimtime="00:00:46.61" lane="6" heatid="5004" />
                <RESULT resultid="1653" eventid="10" swimtime="00:01:40.37" lane="6" heatid="10004" />
                <RESULT resultid="1652" eventid="12" swimtime="00:00:39.39" lane="4" heatid="12008" />
                <RESULT resultid="1651" eventid="17" swimtime="00:01:02.69" lane="4" heatid="17008" />
                <RESULT resultid="1650" eventid="23" swimtime="00:03:13.76" lane="3" heatid="23004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:31.35" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1649" eventid="33" swimtime="00:01:29.73" lane="7" heatid="33009" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="343" birthdate="2014-01-01" gender="F" lastname="Schüller" firstname="Aurelia Ida-Charlotte" license="448124">
              <RESULTS>
                <RESULT resultid="1658" eventid="19" swimtime="00:00:56.68" lane="3" heatid="19012" />
                <RESULT resultid="1657" eventid="25" swimtime="00:00:50.02" lane="3" heatid="25019" />
                <RESULT resultid="1656" eventid="29" swimtime="00:00:40.55" lane="2" heatid="29013" />
                <RESULT resultid="1655" eventid="33" swimtime="00:01:35.82" lane="2" heatid="33005" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="344" birthdate="2014-01-01" gender="F" lastname="Sachse" firstname="Antonia" license="461705">
              <RESULTS>
                <RESULT resultid="1663" eventid="17" swimtime="00:01:05.57" lane="5" heatid="17006" />
                <RESULT resultid="1662" eventid="21" swimtime="00:01:07.86" lane="5" heatid="21008" />
                <RESULT resultid="1661" eventid="25" swimtime="00:00:48.48" lane="3" heatid="25018" />
                <RESULT resultid="1660" eventid="29" swimtime="00:00:43.02" lane="5" heatid="29011" />
                <RESULT resultid="1659" eventid="33" swimtime="00:01:38.44" lane="4" heatid="33002" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="SC Chemnitz von 1892" nation="GER" region="12" code="3353">
          <ATHLETES>
            <ATHLETE athleteid="924" birthdate="2014-01-01" gender="F" lastname="Klimant" firstname="Alexandra" license="448305">
              <RESULTS>
                <RESULT resultid="4326" eventid="17" swimtime="00:01:01.05" lane="6" heatid="17013" />
                <RESULT resultid="4327" eventid="21" swimtime="00:00:57.49" lane="4" heatid="21011" />
                <RESULT resultid="4328" eventid="25" swimtime="00:00:52.08" lane="7" heatid="25017" />
                <RESULT resultid="4329" eventid="29" swimtime="00:00:41.87" lane="8" heatid="29011" />
                <RESULT resultid="4330" eventid="31" swimtime="00:00:56.36" lane="6" heatid="31006" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="925" birthdate="2014-01-01" gender="F" lastname="Pelz" firstname="Alma" license="448311">
              <RESULTS>
                <RESULT resultid="4331" eventid="17" swimtime="00:01:02.89" lane="8" heatid="17011" />
                <RESULT resultid="4332" eventid="21" swimtime="00:01:03.33" lane="3" heatid="21007" />
                <RESULT resultid="4333" eventid="25" swimtime="00:00:48.20" lane="2" heatid="25015" />
                <RESULT resultid="4334" eventid="29" swimtime="00:00:44.78" lane="8" heatid="29013" />
                <RESULT resultid="4335" eventid="31" swimtime="00:01:01.22" lane="4" heatid="31004" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="926" birthdate="2015-01-01" gender="F" lastname="Fehle" firstname="Anni" license="463845">
              <RESULTS>
                <RESULT resultid="4336" eventid="17" swimtime="00:01:00.10" lane="6" heatid="17012" />
                <RESULT resultid="4337" eventid="21" swimtime="00:00:57.64" lane="3" heatid="21008" />
                <RESULT resultid="4338" eventid="25" swimtime="00:00:49.77" lane="5" heatid="25016" />
                <RESULT resultid="4339" eventid="29" swimtime="00:00:43.20" lane="7" heatid="29011" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="927" birthdate="2015-01-01" gender="F" lastname="Kühn" firstname="Antonia" license="458175">
              <RESULTS>
                <RESULT resultid="4340" eventid="19" swimtime="00:00:52.87" lane="1" heatid="19010" />
                <RESULT resultid="4341" eventid="21" swimtime="00:00:56.23" lane="5" heatid="21011" />
                <RESULT resultid="4342" eventid="27" swimtime="00:01:03.07" lane="2" heatid="27011" />
                <RESULT resultid="4343" eventid="29" swimtime="00:00:47.41" lane="1" heatid="29007" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="928" birthdate="2013-01-01" gender="M" lastname="Roßburg" firstname="Ben" license="445426">
              <RESULTS>
                <RESULT resultid="4344" eventid="20" swimtime="00:00:51.38" lane="5" heatid="20012" />
                <RESULT resultid="4345" eventid="24" swimtime="00:03:00.86" lane="7" heatid="24004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:28.12" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="4346" eventid="32" swimtime="00:00:56.62" lane="1" heatid="32004" />
                <RESULT resultid="4347" eventid="36" swimtime="00:01:34.14" lane="7" heatid="36002" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="929" birthdate="2012-01-01" gender="M" lastname="Wendritsch" firstname="Ben" license="437416">
              <RESULTS>
                <RESULT resultid="4348" eventid="18" swimtime="00:00:56.60" lane="1" heatid="18012" />
                <RESULT resultid="4349" eventid="26" swimtime="00:00:42.93" lane="8" heatid="26019" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="930" birthdate="2015-01-01" gender="F" lastname="Mann" firstname="Elisa" license="464000">
              <RESULTS>
                <RESULT resultid="4350" eventid="17" swimtime="00:01:08.11" lane="7" heatid="17006" />
                <RESULT resultid="4351" eventid="21" swimtime="00:01:04.57" lane="4" heatid="21004" />
                <RESULT resultid="4352" eventid="25" swimtime="00:01:04.29" lane="2" heatid="25005" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="931" birthdate="2013-01-01" gender="F" lastname="Maier" firstname="Elli" license="444228">
              <RESULTS>
                <RESULT resultid="4353" eventid="19" swimtime="00:00:56.10" lane="2" heatid="19012" />
                <RESULT resultid="4354" eventid="23" swimtime="00:03:33.71" lane="4" heatid="23001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:42.08" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="4355" eventid="27" swimtime="00:01:02.15" lane="2" heatid="27010" />
                <RESULT resultid="4356" eventid="33" swimtime="00:01:39.17" lane="4" heatid="33003" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="932" birthdate="2013-01-01" gender="F" lastname="Peter" firstname="Emma" license="444231">
              <RESULTS>
                <RESULT resultid="4357" eventid="17" swimtime="00:00:59.65" lane="3" heatid="17014" />
                <RESULT resultid="4358" eventid="25" swimtime="00:00:46.34" lane="3" heatid="25017" />
                <RESULT resultid="4359" eventid="31" swimtime="00:01:01.83" lane="7" heatid="31006" />
                <RESULT resultid="4360" eventid="33" swimtime="00:01:37.71" lane="8" heatid="33005" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="933" birthdate="2014-01-01" gender="F" lastname="Pfeifer" firstname="Feena" license="448306">
              <RESULTS>
                <RESULT resultid="4361" eventid="19" swimtime="00:00:55.90" lane="1" heatid="19008" />
                <RESULT resultid="4362" eventid="21" swimtime="00:01:05.76" lane="6" heatid="21009" />
                <RESULT resultid="4363" eventid="25" swimtime="00:00:48.41" lane="7" heatid="25015" />
                <RESULT resultid="4364" eventid="27" swimtime="00:01:04.90" lane="6" heatid="27009" />
                <RESULT resultid="4365" eventid="31" swimtime="00:01:07.14" lane="7" heatid="31005" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="934" birthdate="2013-01-01" gender="M" lastname="Goebel" firstname="Ferdinand" license="444239">
              <RESULTS>
                <RESULT resultid="4366" eventid="20" swimtime="00:00:43.79" lane="5" heatid="20017" />
                <RESULT resultid="4367" eventid="28" swimtime="00:00:52.80" lane="7" heatid="28008" />
                <RESULT resultid="4368" eventid="32" swimtime="00:00:55.29" lane="3" heatid="32005" />
                <RESULT resultid="4369" eventid="34" swimtime="00:01:27.46" lane="4" heatid="34006" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="935" birthdate="2014-01-01" gender="F" lastname="Kotulla" firstname="Frieda" license="448312">
              <RESULTS>
                <RESULT resultid="4370" eventid="19" swimtime="00:00:58.52" lane="2" heatid="19009" />
                <RESULT resultid="4371" eventid="21" swimtime="00:00:58.23" lane="8" heatid="21013" />
                <RESULT resultid="4372" eventid="25" swimtime="00:00:52.05" lane="7" heatid="25012" />
                <RESULT resultid="4373" eventid="29" swimtime="00:00:42.37" lane="3" heatid="29012" />
                <RESULT resultid="4374" eventid="31" status="DSQ" swimtime="00:01:02.69" lane="8" heatid="31006" comment="Wechselbeinschläge." />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="936" birthdate="2015-01-01" gender="M" lastname="Brandt" firstname="Fritz" license="463996">
              <RESULTS>
                <RESULT resultid="4375" eventid="18" swimtime="00:01:00.54" lane="7" heatid="18010" />
                <RESULT resultid="4376" eventid="20" swimtime="00:00:59.66" lane="8" heatid="20005" />
                <RESULT resultid="4377" eventid="22" swimtime="00:00:56.41" lane="8" heatid="22010" />
                <RESULT resultid="4378" eventid="26" swimtime="00:00:47.57" lane="6" heatid="26008" />
                <RESULT resultid="4379" eventid="30" swimtime="00:00:40.79" lane="4" heatid="30005" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="937" birthdate="2014-01-01" gender="F" lastname="Engmann" firstname="Greta" license="448303">
              <RESULTS>
                <RESULT resultid="4380" eventid="19" swimtime="00:00:51.28" lane="2" heatid="19016" />
                <RESULT resultid="4381" eventid="25" swimtime="00:00:46.87" lane="7" heatid="25020" />
                <RESULT resultid="4382" eventid="29" swimtime="00:00:40.34" lane="3" heatid="29013" />
                <RESULT resultid="4383" eventid="33" swimtime="00:01:33.41" lane="7" heatid="33007" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="938" birthdate="2015-01-01" gender="F" lastname="Rother" firstname="Hannah" license="463855">
              <RESULTS>
                <RESULT resultid="4384" eventid="17" swimtime="00:01:01.86" lane="8" heatid="17010" />
                <RESULT resultid="4385" eventid="21" swimtime="00:01:03.00" lane="4" heatid="21008" />
                <RESULT resultid="4386" eventid="25" swimtime="00:00:54.40" lane="3" heatid="25010" />
                <RESULT resultid="4387" eventid="29" swimtime="00:00:44.12" lane="8" heatid="29008" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="939" birthdate="2011-01-01" gender="F" lastname="Schultze" firstname="Heidi" license="423424">
              <RESULTS>
                <RESULT resultid="4388" eventid="10" swimtime="00:01:29.90" lane="6" heatid="10007" />
                <RESULT resultid="4389" eventid="12" swimtime="00:00:34.80" lane="6" heatid="12012" />
                <RESULT resultid="4390" eventid="23" swimtime="00:02:38.27" lane="3" heatid="23009">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:17.21" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="4391" eventid="25" swimtime="00:00:42.20" lane="1" heatid="25024" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="940" birthdate="2013-01-01" gender="M" lastname="Toth" firstname="Henry" license="444224">
              <RESULTS>
                <RESULT resultid="4392" eventid="22" swimtime="00:00:56.45" lane="1" heatid="22008" />
                <RESULT resultid="4393" eventid="24" swimtime="00:03:00.74" lane="2" heatid="24004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:29.94" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="4394" eventid="34" swimtime="00:01:19.59" lane="5" heatid="34007" />
                <RESULT resultid="4395" eventid="38" status="DSQ" swimtime="00:03:18.96" lane="3" heatid="38001" comment="Bei der 2. Wende wurde die Wende nicht unverzüglich nach Einnahme der Bauchlage ausgeführt.">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:39.04" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="941" birthdate="2015-01-01" gender="M" lastname="Böhm" firstname="Jonas" license="463989">
              <RESULTS>
                <RESULT resultid="4396" eventid="20" swimtime="00:00:55.45" lane="4" heatid="20006" />
                <RESULT resultid="4397" eventid="22" swimtime="00:01:10.49" lane="4" heatid="22004" />
                <RESULT resultid="4398" eventid="28" swimtime="00:01:00.91" lane="5" heatid="28006" />
                <RESULT resultid="4399" eventid="30" swimtime="00:00:46.71" lane="7" heatid="30005" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="942" birthdate="2012-01-01" gender="M" lastname="Li" firstname="Joshua" license="437425">
              <RESULTS>
                <RESULT resultid="4400" eventid="20" swimtime="00:00:42.18" lane="3" heatid="20019" />
                <RESULT resultid="4401" eventid="28" swimtime="00:00:52.92" lane="4" heatid="28008" />
                <RESULT resultid="4402" eventid="32" swimtime="00:00:49.34" lane="5" heatid="32005" />
                <RESULT resultid="4403" eventid="36" swimtime="00:01:26.23" lane="3" heatid="36002" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="943" birthdate="2012-01-01" gender="F" lastname="Herrmann" firstname="Juli" license="437421">
              <RESULTS>
                <RESULT resultid="4404" eventid="17" status="DNS" swimtime="00:00:00.00" lane="2" heatid="17015" />
                <RESULT resultid="4405" eventid="25" status="DNS" swimtime="00:00:00.00" lane="3" heatid="25029" />
                <RESULT resultid="4406" eventid="31" status="DNS" swimtime="00:00:00.00" lane="5" heatid="31007" />
                <RESULT resultid="4407" eventid="37" status="DNS" swimtime="00:00:00.00" lane="6" heatid="37006" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="944" birthdate="2014-01-01" gender="F" lastname="Gottschalk" firstname="Julia" license="448307">
              <RESULTS>
                <RESULT resultid="4408" eventid="19" swimtime="00:00:47.21" lane="6" heatid="19018" />
                <RESULT resultid="4409" eventid="21" swimtime="00:01:05.09" lane="4" heatid="21009" />
                <RESULT resultid="4410" eventid="25" swimtime="00:00:47.89" lane="2" heatid="25019" />
                <RESULT resultid="4411" eventid="27" swimtime="00:01:02.16" lane="1" heatid="27010" />
                <RESULT resultid="4412" eventid="33" swimtime="00:01:36.46" lane="5" heatid="33004" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="945" birthdate="2015-01-01" gender="F" lastname="Hübner" firstname="Julia" license="463859">
              <RESULTS>
                <RESULT resultid="4413" eventid="17" swimtime="00:01:10.38" lane="3" heatid="17004" />
                <RESULT resultid="4414" eventid="21" swimtime="00:01:12.95" lane="5" heatid="21004" />
                <RESULT resultid="4415" eventid="25" status="DSQ" swimtime="00:00:58.41" lane="5" heatid="25005" comment="Anschlag nicht in Rückenlage." />
                <RESULT resultid="4416" eventid="29" swimtime="00:00:57.89" lane="7" heatid="29002" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="946" birthdate="2012-01-01" gender="M" lastname="Barth" firstname="Justus" license="438038">
              <RESULTS>
                <RESULT resultid="4417" eventid="22" swimtime="00:00:47.46" lane="5" heatid="22010" />
                <RESULT resultid="4418" eventid="26" swimtime="00:00:40.17" lane="3" heatid="26020" />
                <RESULT resultid="4419" eventid="34" swimtime="00:01:21.04" lane="7" heatid="34009" />
                <RESULT resultid="4420" eventid="38" swimtime="00:03:14.49" lane="2" heatid="38003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:39.41" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="947" birthdate="2013-01-01" gender="M" lastname="Stark" firstname="Lennart" license="444234">
              <RESULTS>
                <RESULT resultid="4421" eventid="18" swimtime="00:00:58.34" lane="6" heatid="18011" />
                <RESULT resultid="4422" eventid="26" swimtime="00:00:45.53" lane="1" heatid="26015" />
                <RESULT resultid="4423" eventid="32" swimtime="00:00:56.37" lane="6" heatid="32004" />
                <RESULT resultid="4424" eventid="38" swimtime="00:03:28.78" lane="1" heatid="38002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:41.86" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="948" birthdate="2015-01-01" gender="F" lastname="May" firstname="Leonie" license="463853">
              <RESULTS>
                <RESULT resultid="4425" eventid="19" swimtime="00:00:58.51" lane="8" heatid="19008" />
                <RESULT resultid="4426" eventid="27" swimtime="00:01:06.92" lane="3" heatid="27007" />
                <RESULT resultid="4427" eventid="29" swimtime="00:00:52.59" lane="4" heatid="29002" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="949" birthdate="2013-01-01" gender="F" lastname="Hernandez" firstname="Lilly" license="444222">
              <RESULTS>
                <RESULT resultid="4428" eventid="17" swimtime="00:00:56.36" lane="7" heatid="17015" />
                <RESULT resultid="4429" eventid="21" swimtime="00:00:51.93" lane="3" heatid="21014" />
                <RESULT resultid="4430" eventid="31" swimtime="00:00:59.58" lane="8" heatid="31007" />
                <RESULT resultid="4431" eventid="37" status="DSQ" swimtime="00:03:37.77" lane="1" heatid="37002" comment="Bei der 1. Wende wurde die Wende nicht unverzüglich nach Einnahme der Bauchlage ausgeführt.">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:48.77" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="950" birthdate="2014-01-01" gender="F" lastname="Gehre" firstname="Linda" license="448310">
              <RESULTS>
                <RESULT resultid="4432" eventid="19" swimtime="00:00:54.04" lane="1" heatid="19009" />
                <RESULT resultid="4433" eventid="25" swimtime="00:00:50.14" lane="8" heatid="25018" />
                <RESULT resultid="4434" eventid="29" swimtime="00:00:42.09" lane="1" heatid="29012" />
                <RESULT resultid="4435" eventid="33" swimtime="00:01:33.29" lane="8" heatid="33007" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="951" birthdate="2012-01-01" gender="F" lastname="Denner" firstname="Linnea" license="438435">
              <RESULTS>
                <RESULT resultid="4436" eventid="12" swimtime="00:00:31.60" lane="1" heatid="12015" />
                <RESULT resultid="4437" eventid="14" swimtime="00:03:06.22" lane="6" heatid="14007">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:30.99" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="4438" eventid="19" swimtime="00:00:39.97" lane="3" heatid="19025" />
                <RESULT resultid="4439" eventid="23" swimtime="00:02:33.57" lane="3" heatid="23005">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:12.69" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="952" birthdate="2011-01-01" gender="F" lastname="Franke" firstname="Loreley" license="447682">
              <RESULTS>
                <RESULT resultid="4440" eventid="10" swimtime="00:01:21.77" lane="7" heatid="10013" />
                <RESULT resultid="4441" eventid="12" swimtime="00:00:32.91" lane="2" heatid="12013" />
                <RESULT resultid="4442" eventid="19" swimtime="00:00:43.93" lane="5" heatid="19020" />
                <RESULT resultid="4443" eventid="25" swimtime="00:00:38.54" lane="1" heatid="25033" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="953" birthdate="2013-01-01" gender="F" lastname="Tittmann" firstname="Luna" license="444223">
              <RESULTS>
                <RESULT resultid="4444" eventid="19" swimtime="00:00:45.93" lane="8" heatid="19024" />
                <RESULT resultid="4445" eventid="25" swimtime="00:00:42.42" lane="1" heatid="25028" />
                <RESULT resultid="4446" eventid="31" swimtime="00:00:51.50" lane="3" heatid="31007" />
                <RESULT resultid="4447" eventid="35" swimtime="00:01:36.56" lane="7" heatid="35003" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="954" birthdate="2015-01-01" gender="F" lastname="Steuer" firstname="Maria" license="463864">
              <RESULTS>
                <RESULT resultid="4448" eventid="19" swimtime="00:00:57.48" lane="7" heatid="19008" />
                <RESULT resultid="4449" eventid="25" swimtime="00:00:58.21" lane="3" heatid="25004" />
                <RESULT resultid="4450" eventid="27" swimtime="00:01:05.67" lane="4" heatid="27005" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="955" birthdate="2012-01-01" gender="M" lastname="Gehre" firstname="Matti" license="437418">
              <RESULTS>
                <RESULT resultid="4451" eventid="18" swimtime="00:00:54.74" lane="3" heatid="18012" />
                <RESULT resultid="4452" eventid="24" swimtime="00:02:43.35" lane="5" heatid="24007">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:19.60" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="4453" eventid="34" swimtime="00:01:13.83" lane="1" heatid="34012" />
                <RESULT resultid="4454" eventid="38" swimtime="00:03:10.23" lane="2" heatid="38004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:34.74" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="956" birthdate="2013-01-01" gender="F" lastname="Wetzel" firstname="Mia Marie" license="444235">
              <RESULTS>
                <RESULT resultid="4455" eventid="19" swimtime="00:00:45.48" lane="3" heatid="19021" />
                <RESULT resultid="4456" eventid="25" swimtime="00:00:46.08" lane="2" heatid="25027" />
                <RESULT resultid="4457" eventid="27" swimtime="00:00:54.48" lane="5" heatid="27012" />
                <RESULT resultid="4458" eventid="37" swimtime="00:03:17.01" lane="8" heatid="37004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:37.00" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="957" birthdate="2014-01-01" gender="F" lastname="Kult" firstname="Milla" license="448302">
              <RESULTS>
                <RESULT resultid="4459" eventid="17" swimtime="00:01:03.13" lane="4" heatid="17012" />
                <RESULT resultid="4460" eventid="21" status="DSQ" swimtime="00:00:56.07" lane="4" heatid="21012" comment="Das Brett wurde beim Zielanschlag vorn nicht umfasst." />
                <RESULT resultid="4461" eventid="25" swimtime="00:00:48.45" lane="4" heatid="25017" />
                <RESULT resultid="4462" eventid="29" swimtime="00:00:44.49" lane="4" heatid="29007" />
                <RESULT resultid="4463" eventid="31" swimtime="00:01:09.42" lane="3" heatid="31002" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="958" birthdate="2011-01-01" gender="M" lastname="Engmann" firstname="Moritz" license="424576">
              <RESULTS>
                <RESULT resultid="4464" eventid="4" swimtime="00:01:25.33" lane="8" heatid="4010" />
                <RESULT resultid="4465" eventid="6" swimtime="00:00:33.80" lane="5" heatid="6007" />
                <RESULT resultid="4466" eventid="11" swimtime="00:01:19.82" lane="5" heatid="11010" />
                <RESULT resultid="4467" eventid="13" swimtime="00:00:30.78" lane="7" heatid="13014" />
                <RESULT resultid="4468" eventid="20" swimtime="00:00:38.57" lane="7" heatid="20016" />
                <RESULT resultid="4469" eventid="24" swimtime="00:02:28.62" lane="8" heatid="24007">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:11.81" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="959" birthdate="2015-01-01" gender="F" lastname="Hommel" firstname="Naima" license="463852">
              <RESULTS>
                <RESULT resultid="4470" eventid="17" swimtime="00:01:04.20" lane="8" heatid="17008" />
                <RESULT resultid="4471" eventid="21" swimtime="00:01:03.91" lane="8" heatid="21005" />
                <RESULT resultid="4472" eventid="25" swimtime="00:00:59.86" lane="8" heatid="25005" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="960" birthdate="2013-01-01" gender="F" lastname="Günther" firstname="Neele" license="444227">
              <RESULTS>
                <RESULT resultid="4473" eventid="17" swimtime="00:01:07.11" lane="3" heatid="17013" />
                <RESULT resultid="4474" eventid="25" swimtime="00:00:45.57" lane="6" heatid="25020" />
                <RESULT resultid="4475" eventid="33" swimtime="00:01:24.68" lane="6" heatid="33008" />
                <RESULT resultid="4476" eventid="37" swimtime="00:03:24.65" lane="5" heatid="37002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:42.30" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="961" birthdate="2012-01-01" gender="F" lastname="Liebisch" firstname="Nele" license="437420">
              <RESULTS>
                <RESULT resultid="4477" eventid="19" swimtime="00:00:50.90" lane="2" heatid="19017" />
                <RESULT resultid="4478" eventid="23" swimtime="00:02:57.65" lane="3" heatid="23006">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:25.83" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="4479" eventid="25" swimtime="00:00:47.10" lane="8" heatid="25024" />
                <RESULT resultid="4480" eventid="35" swimtime="00:01:45.00" lane="8" heatid="35003" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="962" birthdate="2012-01-01" gender="M" lastname="Naumann" firstname="Nilo" license="444950">
              <RESULTS>
                <RESULT resultid="4481" eventid="22" swimtime="00:00:58.89" lane="5" heatid="22009" />
                <RESULT resultid="4482" eventid="28" swimtime="00:01:03.34" lane="2" heatid="28007" />
                <RESULT resultid="4483" eventid="32" swimtime="00:01:04.29" lane="6" heatid="32005" />
                <RESULT resultid="4484" eventid="34" swimtime="00:01:32.19" lane="5" heatid="34005" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="963" birthdate="2015-01-01" gender="F" lastname="Seidler" firstname="Nina" license="463856">
              <RESULTS>
                <RESULT resultid="4485" eventid="19" swimtime="00:01:03.51" lane="5" heatid="19006" />
                <RESULT resultid="4486" eventid="21" swimtime="00:01:11.70" lane="2" heatid="21004" />
                <RESULT resultid="4487" eventid="27" swimtime="00:01:10.19" lane="8" heatid="27006" />
                <RESULT resultid="4488" eventid="29" swimtime="00:00:56.39" lane="3" heatid="29005" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="964" birthdate="2015-01-01" gender="F" lastname="Sinang" firstname="Nora" license="463857">
              <RESULTS>
                <RESULT resultid="4489" eventid="19" swimtime="00:00:54.89" lane="7" heatid="19012" />
                <RESULT resultid="4490" eventid="25" swimtime="00:00:53.89" lane="3" heatid="25007" />
                <RESULT resultid="4491" eventid="27" swimtime="00:01:01.69" lane="5" heatid="27010" />
                <RESULT resultid="4492" eventid="29" swimtime="00:00:49.40" lane="4" heatid="29005" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="965" birthdate="2015-01-01" gender="M" lastname="Böhm" firstname="Oskar" license="463988">
              <RESULTS>
                <RESULT resultid="4493" eventid="20" swimtime="00:00:59.31" lane="6" heatid="20004" />
                <RESULT resultid="4494" eventid="26" swimtime="00:00:52.83" lane="7" heatid="26007" />
                <RESULT resultid="4495" eventid="28" swimtime="00:01:05.03" lane="4" heatid="28005" />
                <RESULT resultid="4496" eventid="30" swimtime="00:00:46.98" lane="6" heatid="30006" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="966" birthdate="2013-01-01" gender="M" lastname="Fröhlich" firstname="Paul" license="445427">
              <RESULTS>
                <RESULT resultid="4497" eventid="18" swimtime="00:00:54.40" lane="6" heatid="18012" />
                <RESULT resultid="4498" eventid="26" swimtime="00:00:42.52" lane="8" heatid="26017" />
                <RESULT resultid="4499" eventid="28" swimtime="00:00:59.86" lane="4" heatid="28006" />
                <RESULT resultid="4500" eventid="38" swimtime="00:03:13.57" lane="4" heatid="38003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:36.66" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="967" birthdate="2012-01-01" gender="F" lastname="Barthold" firstname="Paula" license="437422">
              <RESULTS>
                <RESULT resultid="4501" eventid="10" swimtime="00:01:29.18" lane="7" heatid="10008" />
                <RESULT resultid="4502" eventid="14" swimtime="00:03:45.99" lane="2" heatid="14004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:49.86" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="4503" eventid="23" swimtime="00:02:56.66" lane="6" heatid="23005">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:25.52" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="4504" eventid="27" status="DNS" swimtime="00:00:00.00" lane="1" heatid="27008" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="968" birthdate="2012-01-01" gender="F" lastname="Drechsel" firstname="Rosalie" license="437426">
              <RESULTS>
                <RESULT resultid="4505" eventid="10" swimtime="00:01:25.13" lane="3" heatid="10011" />
                <RESULT resultid="4506" eventid="14" swimtime="00:03:39.68" lane="5" heatid="14004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:44.66" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="4507" eventid="23" swimtime="00:02:42.01" lane="8" heatid="23008">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:18.79" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="4508" eventid="25" swimtime="00:00:41.06" lane="1" heatid="25030" />
                <RESULT resultid="4509" eventid="37" swimtime="00:03:02.99" lane="1" heatid="37007">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:30.72" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="969" birthdate="2013-01-01" gender="F" lastname="Wild" firstname="Sara" license="444949">
              <RESULTS>
                <RESULT resultid="4510" eventid="21" swimtime="00:00:54.82" lane="6" heatid="21013" />
                <RESULT resultid="4511" eventid="23" swimtime="00:02:54.45" lane="3" heatid="23007">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:25.32" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="4512" eventid="31" swimtime="00:00:52.65" lane="3" heatid="31006" />
                <RESULT resultid="4513" eventid="37" swimtime="00:03:13.02" lane="5" heatid="37003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:35.05" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="970" birthdate="2013-01-01" gender="F" lastname="Keil" firstname="Sophie" license="444232">
              <RESULTS>
                <RESULT resultid="4514" eventid="21" swimtime="00:00:52.33" lane="1" heatid="21014" />
                <RESULT resultid="4515" eventid="23" swimtime="00:02:57.27" lane="2" heatid="23007">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:25.99" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="4516" eventid="33" swimtime="00:01:22.07" lane="6" heatid="33011" />
                <RESULT resultid="4517" eventid="37" swimtime="00:03:27.60" lane="6" heatid="37002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:43.50" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="971" birthdate="2015-01-01" gender="M" lastname="Kechagias" firstname="Thanos" license="464505">
              <RESULTS>
                <RESULT resultid="4518" eventid="20" swimtime="00:00:56.83" lane="3" heatid="20006" />
                <RESULT resultid="4519" eventid="26" swimtime="00:00:53.86" lane="5" heatid="26004" />
                <RESULT resultid="4520" eventid="28" swimtime="00:01:06.38" lane="3" heatid="28004" />
                <RESULT resultid="4521" eventid="30" swimtime="00:00:51.04" lane="5" heatid="30003" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="972" birthdate="2015-01-01" gender="M" lastname="Hecker" firstname="Tom" license="463846">
              <RESULTS>
                <RESULT resultid="4522" eventid="18" swimtime="00:01:02.26" lane="8" heatid="18009" />
                <RESULT resultid="4523" eventid="22" swimtime="00:01:07.38" lane="7" heatid="22004" />
                <RESULT resultid="4524" eventid="26" swimtime="00:00:50.90" lane="8" heatid="26008" />
                <RESULT resultid="4525" eventid="30" swimtime="00:00:47.49" lane="7" heatid="30004" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="973" birthdate="2015-01-01" gender="F" lastname="Lorfing" firstname="Valentina" license="463851">
              <RESULTS>
                <RESULT resultid="4526" eventid="19" swimtime="00:01:00.48" lane="6" heatid="19007" />
                <RESULT resultid="4527" eventid="25" swimtime="00:00:57.44" lane="1" heatid="25008" />
                <RESULT resultid="4528" eventid="27" swimtime="00:01:16.41" lane="5" heatid="27007" />
                <RESULT resultid="4529" eventid="29" swimtime="00:00:52.04" lane="3" heatid="29007" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="SC DHfK Leipzig" nation="GER" region="12" code="3354">
          <ATHLETES>
            <ATHLETE athleteid="142" birthdate="2013-01-01" gender="M" lastname="Valeev" firstname="Zakhar" license="448350">
              <RESULTS>
                <RESULT resultid="760" eventid="20" swimtime="00:00:45.42" lane="6" heatid="20010" />
                <RESULT resultid="759" eventid="26" swimtime="00:00:44.83" lane="6" heatid="26012" />
                <RESULT resultid="758" eventid="34" swimtime="00:01:28.42" lane="6" heatid="34003" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="143" birthdate="2013-01-01" gender="F" lastname="Paschy" firstname="Vivien Elisabeth" license="448339">
              <RESULTS>
                <RESULT resultid="763" eventid="19" swimtime="00:00:52.59" lane="7" heatid="19009" />
                <RESULT resultid="762" eventid="25" swimtime="00:00:46.39" lane="6" heatid="25021" />
                <RESULT resultid="761" eventid="33" swimtime="00:01:33.83" lane="5" heatid="33006" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="144" birthdate="2013-01-01" gender="F" lastname="Lißner" firstname="Phoebe" license="448337">
              <RESULTS>
                <RESULT resultid="766" eventid="19" swimtime="00:00:46.53" lane="2" heatid="19020" />
                <RESULT resultid="765" eventid="25" swimtime="00:00:41.36" lane="1" heatid="25029" />
                <RESULT resultid="764" eventid="35" swimtime="00:01:32.68" lane="5" heatid="35001" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="145" birthdate="2010-01-01" gender="M" lastname="Turich" firstname="Niklas" license="417679">
              <RESULTS>
                <RESULT resultid="774" eventid="2" status="DSQ" swimtime="00:02:45.66" lane="7" heatid="2007" comment="Der Sportler führte nach dem Start mehrere Kraularme aus.">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:18.62" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="773" eventid="4" swimtime="00:01:24.36" lane="4" heatid="4009" />
                <RESULT resultid="772" eventid="13" swimtime="00:00:29.57" lane="3" heatid="13015" />
                <RESULT resultid="771" eventid="15" swimtime="00:03:01.34" lane="5" heatid="15006">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:28.98" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="770" eventid="20" swimtime="00:00:37.61" lane="7" heatid="20017" />
                <RESULT resultid="769" eventid="26" swimtime="00:00:33.65" lane="8" heatid="26024" />
                <RESULT resultid="768" eventid="34" swimtime="00:01:06.84" lane="4" heatid="34013" />
                <RESULT resultid="767" eventid="36" swimtime="00:01:21.70" lane="5" heatid="36002" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="146" birthdate="2011-01-01" gender="M" lastname="Milbach" firstname="Mio Moritz" license="408265">
              <RESULTS>
                <RESULT resultid="777" eventid="20" status="DNS" swimtime="00:00:00.00" lane="3" heatid="20011" />
                <RESULT resultid="776" eventid="26" status="DNS" swimtime="00:00:00.00" lane="7" heatid="26017" />
                <RESULT resultid="775" eventid="34" status="DNS" swimtime="00:00:00.00" lane="1" heatid="34008" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="147" birthdate="2013-01-01" gender="F" lastname="Kirschner" firstname="Luise" license="446727">
              <RESULTS>
                <RESULT resultid="781" eventid="19" swimtime="00:00:51.45" lane="1" heatid="19015" />
                <RESULT resultid="780" eventid="27" swimtime="00:00:59.38" lane="3" heatid="27011" />
                <RESULT resultid="779" eventid="31" swimtime="00:01:08.85" lane="3" heatid="31003" />
                <RESULT resultid="778" eventid="33" swimtime="00:01:39.86" lane="7" heatid="33004" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="148" birthdate="2012-01-01" gender="M" lastname="Luschnitz" firstname="Konstantin Paul" license="444085">
              <RESULTS>
                <RESULT resultid="784" eventid="20" swimtime="00:00:50.41" lane="4" heatid="20012" />
                <RESULT resultid="783" eventid="26" swimtime="00:00:41.57" lane="4" heatid="26017" />
                <RESULT resultid="782" eventid="34" swimtime="00:01:22.73" lane="5" heatid="34006" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="149" birthdate="2013-01-01" gender="F" lastname="Gernegroß" firstname="Elsa" license="446725">
              <RESULTS>
                <RESULT resultid="788" eventid="19" status="DNS" swimtime="00:00:00.00" lane="2" heatid="19011" />
                <RESULT resultid="787" eventid="25" status="DNS" swimtime="00:00:00.00" lane="4" heatid="25014" />
                <RESULT resultid="786" eventid="27" status="DNS" swimtime="00:00:00.00" lane="2" heatid="27009" />
                <RESULT resultid="785" eventid="33" status="DNS" swimtime="00:00:00.00" lane="2" heatid="33003" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="150" birthdate="2010-01-01" gender="M" lastname="Füchsel" firstname="Ben" license="417683">
              <RESULTS>
                <RESULT resultid="796" eventid="2" swimtime="00:02:42.44" lane="5" heatid="2007">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:17.22" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="795" eventid="6" swimtime="00:00:35.13" lane="5" heatid="6008" />
                <RESULT resultid="794" eventid="11" swimtime="00:01:20.97" lane="8" heatid="11011" />
                <RESULT resultid="793" eventid="13" swimtime="00:00:30.69" lane="3" heatid="13014" />
                <RESULT resultid="792" eventid="20" swimtime="00:00:40.84" lane="4" heatid="20019" />
                <RESULT resultid="791" eventid="24" swimtime="00:02:23.96" lane="5" heatid="24008">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:09.38" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="790" eventid="34" swimtime="00:01:07.25" lane="5" heatid="34013" />
                <RESULT resultid="789" eventid="36" swimtime="00:01:19.20" lane="8" heatid="36003" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="151" birthdate="2013-01-01" gender="F" lastname="Möschke" firstname="Antonia" license="448338">
              <RESULTS>
                <RESULT resultid="799" eventid="19" swimtime="00:00:50.96" lane="3" heatid="19016" />
                <RESULT resultid="798" eventid="25" swimtime="00:00:40.07" lane="5" heatid="25028" />
                <RESULT resultid="797" eventid="35" swimtime="00:01:34.63" lane="4" heatid="35001" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="152" birthdate="2014-01-01" gender="F" lastname="Rüger" firstname="Amy" license="446724">
              <RESULTS>
                <RESULT resultid="803" eventid="19" swimtime="00:00:44.79" lane="8" heatid="19021" />
                <RESULT resultid="802" eventid="27" swimtime="00:00:54.12" lane="6" heatid="27012" />
                <RESULT resultid="801" eventid="29" swimtime="00:00:40.69" lane="1" heatid="29013" />
                <RESULT resultid="800" eventid="33" swimtime="00:01:33.78" lane="6" heatid="33004" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="153" birthdate="2012-01-01" gender="F" lastname="Barkawitz" firstname="Lotta" license="426141">
              <RESULTS>
                <RESULT resultid="806" eventid="25" swimtime="00:00:41.23" lane="7" heatid="25031" />
                <RESULT resultid="805" eventid="33" swimtime="00:01:20.97" lane="5" heatid="33010" />
                <RESULT resultid="804" eventid="37" swimtime="00:03:11.90" lane="5" heatid="37004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:32.96" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="154" birthdate="2010-01-01" gender="M" lastname="Belyavskiy" firstname="Alexander" license="426136">
              <RESULTS>
                <RESULT resultid="810" eventid="20" swimtime="00:00:39.93" lane="7" heatid="20019" />
                <RESULT resultid="809" eventid="26" swimtime="00:00:33.23" lane="5" heatid="26023" />
                <RESULT resultid="808" eventid="34" swimtime="00:01:03.56" lane="1" heatid="34015" />
                <RESULT resultid="807" eventid="38" swimtime="00:02:31.69" lane="5" heatid="38005">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:15.18" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="SC DHfK Leipzig Flossenschwimmen" nation="GER" region="20" code="0">
          <ATHLETES>
            <ATHLETE athleteid="313" birthdate="2013-01-01" gender="F" lastname="Amelung" firstname="Tabea" license="0">
              <RESULTS>
                <RESULT resultid="1532" eventid="39" swimtime="00:02:29.82" lane="2" heatid="39002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:14.21" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1531" eventid="41" swimtime="00:00:16.32" lane="8" heatid="41004" />
                <RESULT resultid="1530" eventid="45" swimtime="00:01:08.04" lane="3" heatid="45004" />
                <RESULT resultid="1529" eventid="47" swimtime="00:00:41.76" lane="3" heatid="47002" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="314" birthdate="2008-01-01" gender="F" lastname="Kulchytska" firstname="Polina" license="0">
              <RESULTS>
                <RESULT resultid="1535" eventid="39" swimtime="00:01:53.63" lane="4" heatid="39003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:55.63" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1534" eventid="45" swimtime="00:00:50.80" lane="4" heatid="45006" />
                <RESULT resultid="1533" eventid="47" swimtime="00:00:32.01" lane="4" heatid="47002" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="315" birthdate="2010-01-01" gender="F" lastname="Horenok" firstname="Polina" license="0">
              <RESULTS>
                <RESULT resultid="1538" eventid="41" swimtime="00:00:13.15" lane="3" heatid="41005" />
                <RESULT resultid="1537" eventid="47" swimtime="00:00:34.49" lane="7" heatid="47002" />
                <RESULT resultid="1536" eventid="49" swimtime="00:00:26.11" lane="3" heatid="49005" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="316" birthdate="2012-01-01" gender="M" lastname="Kulchytskyi" firstname="Mykyta" license="0">
              <RESULTS>
                <RESULT resultid="1542" eventid="40" swimtime="00:02:11.90" lane="4" heatid="40002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:03.34" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1541" eventid="42" swimtime="00:00:13.45" lane="2" heatid="42003" />
                <RESULT resultid="1540" eventid="46" swimtime="00:01:01.10" lane="2" heatid="46003" />
                <RESULT resultid="1539" eventid="48" swimtime="00:00:39.24" lane="3" heatid="48001" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="317" birthdate="2011-01-01" gender="F" lastname="Schröter" firstname="Melissa" license="0">
              <RESULTS>
                <RESULT resultid="1546" eventid="39" swimtime="00:02:38.96" lane="4" heatid="39001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:16.96" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1545" eventid="41" swimtime="00:00:16.12" lane="2" heatid="41004" />
                <RESULT resultid="1544" eventid="45" swimtime="00:01:08.67" lane="4" heatid="45003" />
                <RESULT resultid="1543" eventid="47" swimtime="00:00:39.36" lane="2" heatid="47002" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="318" birthdate="2012-01-01" gender="M" lastname="Schnepel" firstname="Marten" license="0">
              <RESULTS>
                <RESULT resultid="1550" eventid="42" swimtime="00:00:15.80" lane="4" heatid="42002" />
                <RESULT resultid="1549" eventid="46" swimtime="00:01:13.68" lane="7" heatid="46002" />
                <RESULT resultid="1548" eventid="48" swimtime="00:00:40.20" lane="7" heatid="48001" />
                <RESULT resultid="1547" eventid="50" swimtime="00:00:32.31" lane="2" heatid="50002" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="319" birthdate="2011-01-01" gender="F" lastname="Reinhardt" firstname="Marla" license="0">
              <RESULTS>
                <RESULT resultid="1554" eventid="41" swimtime="00:00:19.22" lane="8" heatid="41003" />
                <RESULT resultid="1553" eventid="45" swimtime="00:01:22.52" lane="4" heatid="45002" />
                <RESULT resultid="1552" eventid="47" swimtime="00:00:47.31" lane="3" heatid="47001" />
                <RESULT resultid="1551" eventid="49" swimtime="00:00:36.99" lane="1" heatid="49002" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="320" birthdate="2011-01-01" gender="F" lastname="Oesterreich" firstname="Mara" license="0">
              <RESULTS>
                <RESULT resultid="1558" eventid="41" swimtime="00:00:17.33" lane="6" heatid="41002" />
                <RESULT resultid="1557" eventid="45" swimtime="00:01:13.07" lane="6" heatid="45003" />
                <RESULT resultid="1556" eventid="47" swimtime="00:00:49.63" lane="8" heatid="47002" />
                <RESULT resultid="1555" eventid="49" swimtime="00:00:32.21" lane="5" heatid="49002" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="321" birthdate="2008-01-01" gender="F" lastname="Horenok" firstname="Maiia" license="0">
              <RESULTS>
                <RESULT resultid="1560" eventid="41" swimtime="00:00:10.15" lane="4" heatid="41005" />
                <RESULT resultid="1559" eventid="49" swimtime="00:00:20.10" lane="4" heatid="49005" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="322" birthdate="2012-01-01" gender="F" lastname="Kossar" firstname="Lisa" license="0">
              <RESULTS>
                <RESULT resultid="1564" eventid="39" swimtime="00:02:28.91" lane="1" heatid="39002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:12.00" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1563" eventid="41" swimtime="00:00:15.67" lane="7" heatid="41004" />
                <RESULT resultid="1562" eventid="45" swimtime="00:01:06.92" lane="7" heatid="45004" />
                <RESULT resultid="1561" eventid="47" swimtime="00:00:37.70" lane="6" heatid="47002" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="323" birthdate="2013-01-01" gender="F" lastname="Kannenberg" firstname="Lilly" license="0">
              <RESULTS>
                <RESULT resultid="1568" eventid="39" swimtime="00:02:32.25" lane="7" heatid="39002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:11.36" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1567" eventid="41" swimtime="00:00:16.86" lane="6" heatid="41004" />
                <RESULT resultid="1566" eventid="45" swimtime="00:01:07.05" lane="2" heatid="45003" />
                <RESULT resultid="1565" eventid="47" swimtime="00:00:45.31" lane="1" heatid="47002" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="324" birthdate="2008-01-01" gender="M" lastname="Hauk" firstname="Leon" license="0">
              <RESULTS>
                <RESULT resultid="1572" eventid="42" swimtime="00:00:15.03" lane="7" heatid="42003" />
                <RESULT resultid="1571" eventid="46" swimtime="00:01:03.33" lane="4" heatid="46002" />
                <RESULT resultid="1570" eventid="48" swimtime="00:00:36.79" lane="2" heatid="48001" />
                <RESULT resultid="1569" eventid="50" swimtime="00:00:28.05" lane="2" heatid="50003" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="325" birthdate="2012-01-01" gender="F" lastname="Hauk" firstname="Laura" license="0">
              <RESULTS>
                <RESULT resultid="1576" eventid="41" swimtime="00:00:15.94" lane="4" heatid="41002" />
                <RESULT resultid="1575" eventid="45" swimtime="00:01:18.84" lane="5" heatid="45002" />
                <RESULT resultid="1574" eventid="47" swimtime="00:00:40.97" lane="4" heatid="47001" />
                <RESULT resultid="1573" eventid="49" swimtime="00:00:33.13" lane="2" heatid="49002" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="326" birthdate="2008-01-01" gender="F" lastname="Säbisch" firstname="Kyra" license="0">
              <RESULTS>
                <RESULT resultid="1578" eventid="41" swimtime="00:00:10.67" lane="5" heatid="41005" />
                <RESULT resultid="1577" eventid="49" swimtime="00:00:21.43" lane="5" heatid="49005" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="327" birthdate="2011-01-01" gender="F" lastname="Hau" firstname="Hannah" license="0">
              <RESULTS>
                <RESULT resultid="1582" eventid="39" swimtime="00:02:15.78" lane="1" heatid="39003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:02.57" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1581" eventid="41" swimtime="00:00:15.06" lane="3" heatid="41004" />
                <RESULT resultid="1580" eventid="45" swimtime="00:00:59.33" lane="4" heatid="45005" />
                <RESULT resultid="1579" eventid="47" swimtime="00:00:36.25" lane="5" heatid="47002" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="328" birthdate="2014-01-01" gender="F" lastname="Paulmann" firstname="Clara Sophie" license="0">
              <RESULTS>
                <RESULT resultid="1586" eventid="43" swimtime="00:00:19.80" lane="4" heatid="43001" />
                <RESULT resultid="1585" eventid="45" swimtime="00:01:28.60" lane="3" heatid="45002" />
                <RESULT resultid="1584" eventid="47" swimtime="00:00:57.91" lane="6" heatid="47001" />
                <RESULT resultid="1583" eventid="49" swimtime="00:00:39.15" lane="8" heatid="49002" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="329" birthdate="2007-01-01" gender="M" lastname="Schoodt" firstname="Ben Joseph" license="2944">
              <RESULTS>
                <RESULT resultid="1589" eventid="42" swimtime="00:00:09.68" lane="4" heatid="42003" />
                <RESULT resultid="1588" eventid="46" swimtime="00:00:42.18" lane="4" heatid="46003" />
                <RESULT resultid="1587" eventid="48" swimtime="00:00:26.42" lane="4" heatid="48001" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="330" birthdate="2013-01-01" gender="M" lastname="Beyer" firstname="Arved" license="0">
              <RESULTS>
                <RESULT resultid="1592" eventid="42" swimtime="00:00:20.37" lane="6" heatid="42002" />
                <RESULT resultid="1591" eventid="46" status="DNS" swimtime="00:00:00.00" lane="6" heatid="46001" />
                <RESULT resultid="1590" eventid="48" status="DNS" swimtime="00:00:00.00" lane="8" heatid="48001" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="331" birthdate="2008-01-01" gender="M" lastname="Berger" firstname="Alex Michael" license="0">
              <RESULTS>
                <RESULT resultid="1594" eventid="42" swimtime="00:00:10.23" lane="5" heatid="42003" />
                <RESULT resultid="1593" eventid="46" swimtime="00:00:46.33" lane="5" heatid="46003" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="SC Freital" nation="GER" region="12" code="3339">
          <ATHLETES>
            <ATHLETE athleteid="115" birthdate="2009-01-01" gender="F" lastname="Lange" firstname="Alia" license="402584">
              <RESULTS>
                <RESULT resultid="610" eventid="33" swimtime="00:01:02.42" lane="4" heatid="33018" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="116" birthdate="2011-01-01" gender="F" lastname="Jang" firstname="Jule" license="425575">
              <RESULTS>
                <RESULT resultid="611" eventid="3" swimtime="00:01:26.11" lane="2" heatid="3011" />
                <RESULT resultid="612" eventid="23" swimtime="00:02:27.39" lane="6" heatid="23011">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:09.73" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="117" birthdate="2010-01-01" gender="F" lastname="Tetzlaff" firstname="Mina Luisa" license="419267">
              <RESULTS>
                <RESULT resultid="613" eventid="10" swimtime="00:01:16.61" lane="1" heatid="10016" />
                <RESULT resultid="614" eventid="12" swimtime="00:00:29.88" lane="8" heatid="12018" />
                <RESULT resultid="615" eventid="33" swimtime="00:01:05.96" lane="2" heatid="33018" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="SC Plauen 06" nation="GER" region="12" code="6374">
          <ATHLETES>
            <ATHLETE athleteid="1355" birthdate="2013-01-01" gender="M" lastname="Friebel" firstname="Ben" license="449440">
              <RESULTS>
                <RESULT resultid="6266" eventid="18" swimtime="00:01:07.98" lane="3" heatid="18003" />
                <RESULT resultid="6267" eventid="22" swimtime="00:01:11.71" lane="3" heatid="22003" />
                <RESULT resultid="6268" eventid="26" swimtime="00:00:51.13" lane="1" heatid="26009" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1356" birthdate="2012-01-01" gender="M" lastname="Schaller" firstname="Benjamin" license="446153">
              <RESULTS>
                <RESULT resultid="6269" eventid="18" swimtime="00:01:08.35" lane="2" heatid="18002" />
                <RESULT resultid="6270" eventid="20" swimtime="00:00:53.52" lane="3" heatid="20010" />
                <RESULT resultid="6271" eventid="22" swimtime="00:01:04.38" lane="1" heatid="22002" />
                <RESULT resultid="6272" eventid="26" swimtime="00:00:48.09" lane="3" heatid="26013" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1357" birthdate="2009-01-01" gender="F" lastname="Weidhase" firstname="Charlotte" license="382370">
              <RESULTS>
                <RESULT resultid="6273" eventid="1" swimtime="00:02:52.10" lane="7" heatid="1007">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:20.04" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="6274" eventid="5" swimtime="00:00:33.70" lane="1" heatid="5013" />
                <RESULT resultid="6275" eventid="10" swimtime="00:01:19.94" lane="5" heatid="10014" />
                <RESULT resultid="6276" eventid="12" swimtime="00:00:30.91" lane="4" heatid="12016" />
                <RESULT resultid="6363" eventid="33" swimtime="00:01:09.29" lane="8" heatid="33002" />
                <RESULT resultid="6277" eventid="35" swimtime="00:01:19.61" lane="3" heatid="35004" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1358" birthdate="2014-01-01" gender="M" lastname="Drescher" firstname="Eddie" license="461630">
              <RESULTS>
                <RESULT resultid="6278" eventid="18" swimtime="00:01:06.67" lane="8" heatid="18010" />
                <RESULT resultid="6279" eventid="22" swimtime="00:01:05.91" lane="6" heatid="22008" />
                <RESULT resultid="6280" eventid="26" swimtime="00:00:52.66" lane="1" heatid="26010" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1359" birthdate="2011-01-01" gender="F" lastname="Georgi" firstname="Elli" license="445741">
              <RESULTS>
                <RESULT resultid="6281" eventid="3" swimtime="00:01:39.21" lane="2" heatid="3005" />
                <RESULT resultid="6282" eventid="5" swimtime="00:00:41.85" lane="7" heatid="5005" />
                <RESULT resultid="6283" eventid="10" swimtime="00:01:32.59" lane="5" heatid="10007" />
                <RESULT resultid="6284" eventid="12" swimtime="00:00:36.86" lane="8" heatid="12010" />
                <RESULT resultid="6285" eventid="19" swimtime="00:00:44.74" lane="5" heatid="19021" />
                <RESULT resultid="6286" eventid="23" swimtime="00:03:00.78" lane="8" heatid="23005">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:25.82" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="6287" eventid="25" swimtime="00:00:42.21" lane="6" heatid="25027" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1360" birthdate="2014-01-01" gender="F" lastname="Damaske" firstname="Emma" license="464467">
              <RESULTS>
                <RESULT resultid="6288" eventid="17" swimtime="00:01:05.30" lane="6" heatid="17007" />
                <RESULT resultid="6289" eventid="21" swimtime="00:01:06.00" lane="7" heatid="21005" />
                <RESULT resultid="6290" eventid="25" swimtime="00:00:49.85" lane="5" heatid="25011" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1361" birthdate="2012-01-01" gender="M" lastname="Reinel" firstname="Falk" license="443315">
              <RESULTS>
                <RESULT resultid="6291" eventid="2" swimtime="00:03:13.54" lane="8" heatid="2005">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:32.57" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="6292" eventid="6" swimtime="00:00:44.68" lane="8" heatid="6005" />
                <RESULT resultid="6293" eventid="11" swimtime="00:01:31.17" lane="6" heatid="11007" />
                <RESULT resultid="6294" eventid="13" swimtime="00:00:34.27" lane="5" heatid="13010" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1362" birthdate="2015-01-01" gender="F" lastname="Schuch" firstname="Finya" license="465816">
              <RESULTS>
                <RESULT resultid="6295" eventid="19" swimtime="00:00:52.86" lane="5" heatid="19011" />
                <RESULT resultid="6296" eventid="21" swimtime="00:00:59.01" lane="7" heatid="21012" />
                <RESULT resultid="6297" eventid="25" swimtime="00:00:48.13" lane="8" heatid="25016" />
                <RESULT resultid="6298" eventid="27" swimtime="00:00:56.48" lane="7" heatid="27012" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1363" birthdate="2012-01-01" gender="M" lastname="Arab" firstname="Hanif Sheikh" license="470911">
              <RESULTS>
                <RESULT resultid="6299" eventid="18" swimtime="00:01:19.89" lane="1" heatid="18002" />
                <RESULT resultid="6300" eventid="22" swimtime="00:01:11.28" lane="6" heatid="22001" />
                <RESULT resultid="6301" eventid="26" swimtime="00:01:00.54" lane="5" heatid="26003" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1364" birthdate="2012-01-01" gender="F" lastname="Fricke" firstname="Helene Hanna" license="443316">
              <RESULTS>
                <RESULT resultid="6302" eventid="17" swimtime="00:01:11.98" lane="2" heatid="17007" />
                <RESULT resultid="6303" eventid="19" swimtime="00:00:52.91" lane="8" heatid="19014" />
                <RESULT resultid="6304" eventid="25" swimtime="00:00:46.36" lane="6" heatid="25019" />
                <RESULT resultid="6305" eventid="27" swimtime="00:01:03.48" lane="8" heatid="27009" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1365" birthdate="2007-01-01" gender="M" lastname="Dressel" firstname="Justin" license="369306">
              <RESULTS>
                <RESULT resultid="6306" eventid="20" swimtime="00:00:36.94" lane="5" heatid="20021" />
                <RESULT resultid="6307" eventid="24" swimtime="00:02:25.45" lane="8" heatid="24009">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:09.65" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="6308" eventid="26" swimtime="00:00:33.33" lane="1" heatid="26024" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1366" birthdate="2011-01-01" gender="M" lastname="Pulz" firstname="Lennox" license="423595">
              <RESULTS>
                <RESULT resultid="6309" eventid="20" swimtime="00:00:49.90" lane="2" heatid="20012" />
                <RESULT resultid="6310" eventid="24" swimtime="00:02:52.30" lane="3" heatid="24004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:25.60" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="6311" eventid="26" swimtime="00:00:45.63" lane="6" heatid="26016" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1367" birthdate="2013-01-01" gender="M" lastname="Pulz" firstname="Liam" license="444209">
              <RESULTS>
                <RESULT resultid="6312" eventid="18" swimtime="00:01:06.73" lane="1" heatid="18004" />
                <RESULT resultid="6313" eventid="20" swimtime="00:00:56.33" lane="4" heatid="20009" />
                <RESULT resultid="6314" eventid="26" swimtime="00:00:51.68" lane="3" heatid="26010" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1368" birthdate="2012-01-01" gender="F" lastname="Uhlig" firstname="Marielle" license="439077">
              <RESULTS>
                <RESULT resultid="6315" eventid="3" swimtime="00:01:37.41" lane="7" heatid="3008" />
                <RESULT resultid="6316" eventid="5" swimtime="00:00:42.76" lane="3" heatid="5005" />
                <RESULT resultid="6317" eventid="10" swimtime="00:01:33.24" lane="6" heatid="10008" />
                <RESULT resultid="6318" eventid="14" swimtime="00:03:32.31" lane="2" heatid="14005">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:44.98" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1369" birthdate="2014-01-01" gender="F" lastname="Feig" firstname="Merle" license="449308">
              <RESULTS>
                <RESULT resultid="6319" eventid="17" status="DNS" swimtime="00:00:00.00" lane="5" heatid="17005" />
                <RESULT resultid="6320" eventid="19" status="DNS" swimtime="00:00:00.00" lane="6" heatid="19010" />
                <RESULT resultid="6321" eventid="25" status="DNS" swimtime="00:00:00.00" lane="3" heatid="25014" />
                <RESULT resultid="6322" eventid="27" status="DNS" swimtime="00:00:00.00" lane="2" heatid="27007" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1370" birthdate="2013-01-01" gender="F" lastname="Gieschke" firstname="Mia" license="444210">
              <RESULTS>
                <RESULT resultid="6323" eventid="17" status="DSQ" swimtime="00:01:11.16" lane="7" heatid="17003" comment="Start vor dem Startsignal." />
                <RESULT resultid="6324" eventid="19" swimtime="00:00:57.36" lane="6" heatid="19008" />
                <RESULT resultid="6325" eventid="25" swimtime="00:00:53.85" lane="7" heatid="25013" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1371" birthdate="2010-01-01" gender="M" lastname="Schreyer" firstname="Miron" license="418771">
              <RESULTS>
                <RESULT resultid="6326" eventid="2" swimtime="00:03:09.33" lane="7" heatid="2005">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:31.78" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="6327" eventid="6" swimtime="00:00:42.53" lane="1" heatid="6006" />
                <RESULT resultid="6328" eventid="11" swimtime="00:01:32.81" lane="1" heatid="11008" />
                <RESULT resultid="6329" eventid="13" swimtime="00:00:34.99" lane="8" heatid="13011" />
                <RESULT resultid="6330" eventid="20" swimtime="00:00:50.69" lane="8" heatid="20013" />
                <RESULT resultid="6331" eventid="24" swimtime="00:02:46.69" lane="1" heatid="24008">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:19.37" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="6332" eventid="26" swimtime="00:00:42.59" lane="6" heatid="26018" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1372" birthdate="2012-01-01" gender="F" lastname="Pöhlmann" firstname="Paula" license="439075">
              <RESULTS>
                <RESULT resultid="6333" eventid="17" swimtime="00:00:55.06" lane="1" heatid="17010" />
                <RESULT resultid="6334" eventid="21" swimtime="00:00:54.07" lane="7" heatid="21010" />
                <RESULT resultid="6335" eventid="25" swimtime="00:00:39.85" lane="4" heatid="25028" />
                <RESULT resultid="6336" eventid="27" swimtime="00:01:07.79" lane="5" heatid="27005" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1373" birthdate="2012-01-01" gender="F" lastname="Breuer" firstname="Pia" license="458559">
              <RESULTS>
                <RESULT resultid="6337" eventid="10" swimtime="00:01:40.56" lane="5" heatid="10004" />
                <RESULT resultid="6338" eventid="12" swimtime="00:00:40.09" lane="3" heatid="12005" />
                <RESULT resultid="6339" eventid="17" swimtime="00:00:55.96" lane="4" heatid="17015" />
                <RESULT resultid="6340" eventid="21" swimtime="00:00:59.76" lane="5" heatid="21014" />
                <RESULT resultid="6341" eventid="25" swimtime="00:00:47.66" lane="1" heatid="25018" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1374" birthdate="2014-01-01" gender="M" lastname="Schaller" firstname="Sebastian" license="449305">
              <RESULTS>
                <RESULT resultid="6342" eventid="20" swimtime="00:01:05.51" lane="1" heatid="20005" />
                <RESULT resultid="6343" eventid="26" swimtime="00:00:54.94" lane="2" heatid="26007" />
                <RESULT resultid="6344" eventid="28" swimtime="00:01:10.14" lane="5" heatid="28004" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1375" birthdate="2012-01-01" gender="F" lastname="Rössel" firstname="Stella" license="439076">
              <RESULTS>
                <RESULT resultid="6345" eventid="10" swimtime="00:01:30.69" lane="6" heatid="10003" />
                <RESULT resultid="6346" eventid="14" swimtime="00:03:25.59" lane="6" heatid="14004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:37.73" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="6347" eventid="19" swimtime="00:00:42.41" lane="8" heatid="19025" />
                <RESULT resultid="6348" eventid="23" swimtime="00:02:49.75" lane="6" heatid="23003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:19.72" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1376" birthdate="2006-01-01" gender="F" lastname="Gruber" firstname="Tessa" license="353903">
              <RESULTS>
                <RESULT resultid="6349" eventid="1" swimtime="00:02:32.57" lane="4" heatid="1007">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:15.29" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="6350" eventid="5" swimtime="00:00:29.44" lane="7" heatid="5014" />
                <RESULT resultid="6351" eventid="10" swimtime="00:01:15.88" lane="6" heatid="10014" />
                <RESULT resultid="6352" eventid="12" swimtime="00:00:27.86" lane="3" heatid="12018" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1377" birthdate="2014-01-01" gender="M" lastname="Wilde" firstname="Vasco" license="454060">
              <RESULTS>
                <RESULT resultid="6353" eventid="18" swimtime="00:01:14.95" lane="6" heatid="18002" />
                <RESULT resultid="6354" eventid="20" swimtime="00:01:01.96" lane="3" heatid="20003" />
                <RESULT resultid="6355" eventid="26" swimtime="00:00:59.74" lane="8" heatid="26005" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1378" birthdate="2014-01-01" gender="M" lastname="Reimann" firstname="Viktor" license="449310">
              <RESULTS>
                <RESULT resultid="6356" eventid="18" swimtime="00:01:06.89" lane="1" heatid="18006" />
                <RESULT resultid="6357" eventid="22" swimtime="00:01:11.11" lane="6" heatid="22003" />
                <RESULT resultid="6358" eventid="26" swimtime="00:00:51.47" lane="6" heatid="26010" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="SC Poseidon Radebeul" nation="GER" region="12" code="3355">
          <ATHLETES>
            <ATHLETE athleteid="1002" birthdate="2015-01-01" gender="M" lastname="Raum" firstname="Fridolin" license="465748">
              <RESULTS>
                <RESULT resultid="4665" eventid="18" swimtime="00:01:06.68" lane="4" heatid="18008" />
                <RESULT resultid="4666" eventid="22" swimtime="00:01:09.43" lane="4" heatid="22006" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1003" birthdate="2015-01-01" gender="F" lastname="Härtwig" firstname="Frieda" license="465755">
              <RESULTS>
                <RESULT resultid="4667" eventid="17" swimtime="00:01:11.20" lane="4" heatid="17011" />
                <RESULT resultid="4668" eventid="21" swimtime="00:01:13.40" lane="3" heatid="21009" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1004" birthdate="2015-01-01" gender="F" lastname="Eichner" firstname="Jette" license="465750">
              <RESULTS>
                <RESULT resultid="4669" eventid="17" status="DNS" swimtime="00:00:00.00" lane="7" heatid="17010" />
                <RESULT resultid="4670" eventid="21" status="DNS" swimtime="00:00:00.00" lane="4" heatid="21007" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1005" birthdate="2007-01-01" gender="F" lastname="Selle" firstname="Marie Elisabeth" license="348768">
              <RESULTS>
                <RESULT resultid="4671" eventid="1" swimtime="00:02:29.03" lane="5" heatid="1007">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:10.80" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="4672" eventid="5" swimtime="00:00:30.30" lane="3" heatid="5014" />
                <RESULT resultid="4673" eventid="10" swimtime="00:01:11.24" lane="5" heatid="10016" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1006" birthdate="2015-01-01" gender="M" lastname="Richter" firstname="Maximilian" license="465958">
              <RESULTS>
                <RESULT resultid="4674" eventid="18" swimtime="00:01:01.99" lane="6" heatid="18007" />
                <RESULT resultid="4675" eventid="20" swimtime="00:00:56.33" lane="3" heatid="20008" />
                <RESULT resultid="4676" eventid="22" swimtime="00:01:07.02" lane="4" heatid="22007" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="SC Riesa" nation="GER" region="12" code="3356">
          <ATHLETES>
            <ATHLETE athleteid="859" birthdate="2010-01-01" gender="M" lastname="Koppe" firstname="Antonio" license="394881">
              <RESULTS>
                <RESULT resultid="4020" eventid="2" swimtime="00:03:09.51" lane="5" heatid="2005">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:23.47" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="4021" eventid="6" swimtime="00:00:35.83" lane="8" heatid="6009" />
                <RESULT resultid="4022" eventid="11" swimtime="00:01:22.17" lane="1" heatid="11011" />
                <RESULT resultid="4023" eventid="13" swimtime="00:00:31.19" lane="5" heatid="13014" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="860" birthdate="2014-01-01" gender="M" lastname="Treptow" firstname="Charlie" license="449100">
              <RESULTS>
                <RESULT resultid="4024" eventid="20" swimtime="00:00:52.83" lane="6" heatid="20009" />
                <RESULT resultid="4025" eventid="26" status="DNS" swimtime="00:00:00.00" lane="3" heatid="26012" />
                <RESULT resultid="4026" eventid="30" status="DNS" swimtime="00:00:00.00" lane="7" heatid="30008" />
                <RESULT resultid="4027" eventid="34" status="DNS" swimtime="00:00:00.00" lane="3" heatid="34002" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="861" birthdate="2011-01-01" gender="F" lastname="Kretzschmar" firstname="Edda-Fränze" license="418095">
              <RESULTS>
                <RESULT resultid="4028" eventid="1" swimtime="00:03:16.93" lane="6" heatid="1004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:35.87" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="4029" eventid="3" swimtime="00:01:37.05" lane="7" heatid="3010" />
                <RESULT resultid="4030" eventid="12" swimtime="00:00:34.30" lane="4" heatid="12012" />
                <RESULT resultid="4031" eventid="14" swimtime="00:03:28.40" lane="2" heatid="14006">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:40.79" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="862" birthdate="2014-01-01" gender="M" lastname="Brade" firstname="Felix" license="449227">
              <RESULTS>
                <RESULT resultid="4032" eventid="20" swimtime="00:00:56.15" lane="8" heatid="20008" />
                <RESULT resultid="4033" eventid="22" swimtime="00:01:12.77" lane="8" heatid="22005" />
                <RESULT resultid="4034" eventid="26" swimtime="00:00:48.79" lane="4" heatid="26011" />
                <RESULT resultid="4035" eventid="30" swimtime="00:00:43.55" lane="4" heatid="30007" />
                <RESULT resultid="4036" eventid="32" swimtime="00:01:06.73" lane="5" heatid="32003" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="863" birthdate="2013-01-01" gender="M" lastname="Thomas" firstname="Florin" license="437788">
              <RESULTS>
                <RESULT resultid="4037" eventid="2" status="DSQ" swimtime="00:03:18.25" lane="2" heatid="2004" comment="Teilstrecke Rücken nicht in Rückenlage beendet.">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:42.28" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="4038" eventid="4" swimtime="00:01:40.68" lane="2" heatid="4007" />
                <RESULT resultid="4039" eventid="13" swimtime="00:00:35.83" lane="2" heatid="13008" />
                <RESULT resultid="4040" eventid="15" swimtime="00:03:31.23" lane="2" heatid="15003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:43.53" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="4041" eventid="20" swimtime="00:00:44.30" lane="2" heatid="20015" />
                <RESULT resultid="4042" eventid="24" swimtime="00:03:01.61" lane="8" heatid="24005">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:27.72" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="4043" eventid="32" swimtime="00:01:08.66" lane="2" heatid="32002" />
                <RESULT resultid="4044" eventid="34" swimtime="00:01:22.53" lane="4" heatid="34007" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="864" birthdate="2014-01-01" gender="M" lastname="Lehmann" firstname="Jonas" license="449099">
              <RESULTS>
                <RESULT resultid="4045" eventid="20" swimtime="00:00:53.36" lane="2" heatid="20008" />
                <RESULT resultid="4046" eventid="22" swimtime="00:01:03.58" lane="3" heatid="22007" />
                <RESULT resultid="4047" eventid="26" swimtime="00:00:48.91" lane="7" heatid="26012" />
                <RESULT resultid="4048" eventid="30" swimtime="00:00:43.35" lane="8" heatid="30008" />
                <RESULT resultid="4049" eventid="34" swimtime="00:01:37.52" lane="2" heatid="34002" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="865" birthdate="2013-01-01" gender="M" lastname="Schäfer" firstname="Jonas" license="449096">
              <RESULTS>
                <RESULT resultid="4050" eventid="6" swimtime="00:00:44.07" lane="1" heatid="6004" />
                <RESULT resultid="4051" eventid="13" swimtime="00:00:36.82" lane="2" heatid="13006" />
                <RESULT resultid="4052" eventid="20" swimtime="00:00:49.54" lane="2" heatid="20013" />
                <RESULT resultid="4053" eventid="26" swimtime="00:00:45.44" lane="7" heatid="26015" />
                <RESULT resultid="4054" eventid="34" swimtime="00:01:22.02" lane="8" heatid="34007" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="866" birthdate="2015-01-01" gender="F" lastname="Cienk" firstname="Klara" license="474171">
              <RESULTS>
                <RESULT resultid="4055" eventid="19" swimtime="00:01:11.58" lane="1" heatid="19001" />
                <RESULT resultid="4056" eventid="21" swimtime="00:01:13.44" lane="3" heatid="21001" />
                <RESULT resultid="4057" eventid="25" swimtime="00:01:08.86" lane="5" heatid="25001" />
                <RESULT resultid="4058" eventid="27" swimtime="00:01:17.62" lane="1" heatid="27002" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="867" birthdate="2010-01-01" gender="F" lastname="Loßner" firstname="Laura" license="376544">
              <RESULTS>
                <RESULT resultid="4059" eventid="1" swimtime="00:03:02.64" lane="8" heatid="1005">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:25.77" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="4060" eventid="5" swimtime="00:00:35.28" lane="4" heatid="5011" />
                <RESULT resultid="4061" eventid="10" swimtime="00:01:27.04" lane="4" heatid="10013" />
                <RESULT resultid="4062" eventid="12" swimtime="00:00:31.94" lane="1" heatid="12017" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="868" birthdate="2012-01-01" gender="M" lastname="Dentel" firstname="Luca" license="422953">
              <RESULTS>
                <RESULT resultid="4063" eventid="2" swimtime="00:03:29.20" lane="1" heatid="2005">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:40.27" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="4064" eventid="4" swimtime="00:01:47.94" lane="5" heatid="4005" />
                <RESULT resultid="4065" eventid="11" swimtime="00:01:39.85" lane="1" heatid="11007" />
                <RESULT resultid="4066" eventid="13" swimtime="00:00:34.15" lane="3" heatid="13010" />
                <RESULT resultid="4067" eventid="20" swimtime="00:00:46.95" lane="2" heatid="20016" />
                <RESULT resultid="4068" eventid="24" swimtime="00:02:59.09" lane="8" heatid="24006">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:27.01" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="4069" eventid="26" swimtime="00:00:42.34" lane="6" heatid="26019" />
                <RESULT resultid="4070" eventid="34" swimtime="00:01:20.27" lane="6" heatid="34010" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="869" birthdate="2010-01-01" gender="F" lastname="Baumgart" firstname="Maria" license="394747">
              <RESULTS>
                <RESULT resultid="4071" eventid="3" status="DNS" swimtime="00:00:00.00" lane="2" heatid="3010" />
                <RESULT resultid="4072" eventid="5" status="DNS" swimtime="00:00:00.00" lane="4" heatid="5006" />
                <RESULT resultid="4073" eventid="12" status="DNS" swimtime="00:00:00.00" lane="3" heatid="12013" />
                <RESULT resultid="4074" eventid="14" status="DNS" swimtime="00:00:00.00" lane="8" heatid="14006" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="870" birthdate="2010-01-01" gender="M" lastname="Brade" firstname="Maximilian" license="394880">
              <RESULTS>
                <RESULT resultid="4075" eventid="2" swimtime="00:03:12.11" lane="4" heatid="2005">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:33.16" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="4076" eventid="11" swimtime="00:01:30.56" lane="1" heatid="11009" />
                <RESULT resultid="4077" eventid="13" swimtime="00:00:36.28" lane="2" heatid="13009" />
                <RESULT resultid="4078" eventid="15" swimtime="00:03:51.04" lane="8" heatid="15004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:55.73" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="871" birthdate="2015-01-01" gender="M" lastname="Zschiegner" firstname="Maximilian" license="457362">
              <RESULTS>
                <RESULT resultid="4079" eventid="18" swimtime="00:01:11.04" lane="5" heatid="18001" />
                <RESULT resultid="4080" eventid="20" swimtime="00:01:07.31" lane="1" heatid="20001" />
                <RESULT resultid="4081" eventid="26" swimtime="00:01:00.61" lane="3" heatid="26001" />
                <RESULT resultid="4082" eventid="28" swimtime="00:01:10.60" lane="4" heatid="28001" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="872" birthdate="2014-01-01" gender="F" lastname="Brade" firstname="Melinda" license="449102">
              <RESULTS>
                <RESULT resultid="4083" eventid="19" swimtime="00:00:57.03" lane="3" heatid="19009" />
                <RESULT resultid="4084" eventid="25" swimtime="00:00:54.56" lane="5" heatid="25012" />
                <RESULT resultid="4085" eventid="29" swimtime="00:00:46.56" lane="2" heatid="29011" />
                <RESULT resultid="4086" eventid="31" swimtime="00:01:12.16" lane="1" heatid="31003" />
                <RESULT resultid="4087" eventid="33" swimtime="00:01:45.11" lane="5" heatid="33003" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="873" birthdate="2015-01-01" gender="F" lastname="Lorenz" firstname="Nele Charlotte" license="457373">
              <RESULTS>
                <RESULT resultid="4088" eventid="17" swimtime="00:01:17.72" lane="1" heatid="17001" />
                <RESULT resultid="4089" eventid="21" swimtime="00:01:10.48" lane="7" heatid="21002" />
                <RESULT resultid="4090" eventid="25" swimtime="00:00:57.55" lane="8" heatid="25007" />
                <RESULT resultid="4091" eventid="27" swimtime="00:01:09.87" lane="1" heatid="27007" />
                <RESULT resultid="4092" eventid="29" swimtime="00:01:03.90" lane="1" heatid="29005" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="874" birthdate="2014-01-01" gender="F" lastname="Sander" firstname="Nicole" license="449231">
              <RESULTS>
                <RESULT resultid="4093" eventid="19" swimtime="00:01:03.67" lane="8" heatid="19006" />
                <RESULT resultid="4094" eventid="25" swimtime="00:00:58.07" lane="6" heatid="25011" />
                <RESULT resultid="4095" eventid="29" swimtime="00:00:49.41" lane="1" heatid="29009" />
                <RESULT resultid="4096" eventid="33" swimtime="00:02:01.32" lane="7" heatid="33002" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="875" birthdate="2013-01-01" gender="M" lastname="Mühlmann" firstname="Ole" license="446953">
              <RESULTS>
                <RESULT resultid="4097" eventid="4" swimtime="00:01:47.93" lane="4" heatid="4004" />
                <RESULT resultid="4098" eventid="13" swimtime="00:00:38.21" lane="5" heatid="13003" />
                <RESULT resultid="4099" eventid="15" swimtime="00:03:54.42" lane="3" heatid="15002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:56.13" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="4100" eventid="20" swimtime="00:00:48.12" lane="3" heatid="20012" />
                <RESULT resultid="4101" eventid="26" swimtime="00:00:43.63" lane="3" heatid="26011" />
                <RESULT resultid="4102" eventid="34" swimtime="00:01:29.91" lane="2" heatid="34004" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="876" birthdate="2008-01-01" gender="M" lastname="Müller" firstname="Stefan" license="384774">
              <RESULTS>
                <RESULT resultid="4103" eventid="4" swimtime="00:01:31.17" lane="6" heatid="4010" />
                <RESULT resultid="4104" eventid="6" swimtime="00:00:29.74" lane="7" heatid="6011" />
                <RESULT resultid="4105" eventid="13" swimtime="00:00:27.01" lane="6" heatid="13018" />
                <RESULT resultid="4106" eventid="15" swimtime="00:03:31.57" lane="5" heatid="15007">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:38.90" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="877" birthdate="2011-01-01" gender="F" lastname="Große" firstname="Viktoria" license="418106">
              <RESULTS>
                <RESULT resultid="4107" eventid="3" swimtime="00:01:43.29" lane="4" heatid="3006" />
                <RESULT resultid="4108" eventid="10" swimtime="00:01:49.08" lane="3" heatid="10004" />
                <RESULT resultid="4109" eventid="12" swimtime="00:00:39.03" lane="5" heatid="12005" />
                <RESULT resultid="4110" eventid="14" swimtime="00:03:48.48" lane="6" heatid="14003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:53.47" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="SC Riesa (TC)" nation="GER" region="20" code="154149">
          <ATHLETES>
            <ATHLETE athleteid="5" birthdate="2011-01-01" gender="F" lastname="Hönisch" firstname="Ida" license="0">
              <RESULTS>
                <RESULT resultid="25" eventid="39" swimtime="00:02:24.29" lane="3" heatid="39002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:08.61" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="26" eventid="41" swimtime="00:00:15.01" lane="6" heatid="41003" />
                <RESULT resultid="27" eventid="45" swimtime="00:01:03.64" lane="5" heatid="45005" />
                <RESULT resultid="28" eventid="49" swimtime="00:00:28.25" lane="6" heatid="49004" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="6" birthdate="2010-01-01" gender="F" lastname="Berger" firstname="Lene" license="0">
              <RESULTS>
                <RESULT resultid="29" eventid="39" swimtime="00:02:15.07" lane="2" heatid="39003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:01.91" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="30" eventid="41" swimtime="00:00:14.22" lane="4" heatid="41004" />
                <RESULT resultid="31" eventid="45" swimtime="00:00:59.29" lane="2" heatid="45006" />
                <RESULT resultid="32" eventid="49" swimtime="00:00:26.66" lane="1" heatid="49005" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="7" birthdate="2014-01-01" gender="F" lastname="Näther" firstname="Mathilde" license="0">
              <RESULTS>
                <RESULT resultid="33" eventid="39" swimtime="00:03:38.31" lane="7" heatid="39001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:39.74" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="34" eventid="43" swimtime="00:00:21.65" lane="3" heatid="43001" />
                <RESULT resultid="35" eventid="45" swimtime="00:01:45.19" lane="7" heatid="45002" />
                <RESULT resultid="36" eventid="49" swimtime="00:00:44.14" lane="6" heatid="49001" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="8" birthdate="2014-01-01" gender="M" lastname="Fleck" firstname="Maximilian" license="0">
              <RESULTS>
                <RESULT resultid="37" eventid="40" swimtime="00:04:12.15" lane="2" heatid="40001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:02:04.28" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="38" eventid="44" swimtime="00:00:30.11" lane="3" heatid="44001" />
                <RESULT resultid="39" eventid="46" swimtime="00:02:04.98" lane="1" heatid="46001" />
                <RESULT resultid="40" eventid="50" swimtime="00:00:57.62" lane="3" heatid="50001" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="9" birthdate="2015-01-01" gender="F" lastname="Sorgalla" firstname="Miriam" license="0">
              <RESULTS>
                <RESULT resultid="41" eventid="39" swimtime="00:03:20.65" lane="2" heatid="39001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:32.49" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="42" eventid="43" swimtime="00:00:21.87" lane="5" heatid="43001" />
                <RESULT resultid="43" eventid="45" swimtime="00:01:36.43" lane="6" heatid="45002" />
                <RESULT resultid="44" eventid="49" swimtime="00:00:42.78" lane="3" heatid="49001" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="10" birthdate="2014-01-01" gender="M" lastname="vom Hoff" firstname="Neo" license="0">
              <RESULTS>
                <RESULT resultid="45" eventid="40" swimtime="00:03:54.87" lane="7" heatid="40001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:52.06" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="46" eventid="44" swimtime="00:00:22.87" lane="5" heatid="44001" />
                <RESULT resultid="47" eventid="46" swimtime="00:01:54.17" lane="7" heatid="46001" />
                <RESULT resultid="48" eventid="50" swimtime="00:00:48.69" lane="5" heatid="50001" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="SSG Leipzig e.V." nation="GER" region="12" code="6466">
          <ATHLETES>
            <ATHLETE athleteid="25" birthdate="2011-01-01" gender="M" lastname="Schmidt" firstname="Arno" license="426924">
              <RESULTS>
                <RESULT resultid="113" eventid="2" swimtime="00:02:54.07" lane="4" heatid="2006">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:20.85" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="114" eventid="6" swimtime="00:00:33.07" lane="6" heatid="6009" />
                <RESULT resultid="115" eventid="11" swimtime="00:01:19.91" lane="3" heatid="11011" />
                <RESULT resultid="116" eventid="13" swimtime="00:00:32.31" lane="2" heatid="13013" />
                <RESULT resultid="117" eventid="20" swimtime="00:00:40.65" lane="5" heatid="20018" />
                <RESULT resultid="118" eventid="26" swimtime="00:00:36.72" lane="6" heatid="26022" />
                <RESULT resultid="119" eventid="34" swimtime="00:01:10.28" lane="4" heatid="34012" />
                <RESULT resultid="120" eventid="38" swimtime="00:02:49.21" lane="7" heatid="38005">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:23.31" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="26" birthdate="2012-01-01" gender="M" lastname="Severyuk" firstname="Daniel" license="440973">
              <RESULTS>
                <RESULT resultid="121" eventid="2" swimtime="00:02:45.72" lane="6" heatid="2007">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:17.80" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="122" eventid="6" swimtime="00:00:31.94" lane="5" heatid="6009" />
                <RESULT resultid="123" eventid="11" swimtime="00:01:17.63" lane="7" heatid="11011" />
                <RESULT resultid="124" eventid="13" swimtime="00:00:30.10" lane="4" heatid="13015" />
                <RESULT resultid="125" eventid="18" swimtime="00:00:44.36" lane="4" heatid="18012" />
                <RESULT resultid="126" eventid="24" swimtime="00:02:26.89" lane="1" heatid="24009">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:11.80" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="127" eventid="34" swimtime="00:01:07.06" lane="3" heatid="34013" />
                <RESULT resultid="128" eventid="38" swimtime="00:02:43.95" lane="8" heatid="38005">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:21.34" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="27" birthdate="2011-01-01" gender="F" lastname="Milbach" firstname="Fanny Madita" license="408264">
              <RESULTS>
                <RESULT resultid="129" eventid="3" swimtime="00:01:26.47" lane="1" heatid="3011" />
                <RESULT resultid="130" eventid="5" swimtime="00:00:33.61" lane="3" heatid="5012" />
                <RESULT resultid="131" eventid="12" swimtime="00:00:31.17" lane="3" heatid="12016" />
                <RESULT resultid="132" eventid="14" swimtime="00:03:08.17" lane="3" heatid="14007">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:30.26" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="133" eventid="19" swimtime="00:00:39.38" lane="3" heatid="19026" />
                <RESULT resultid="134" eventid="25" swimtime="00:00:34.40" lane="3" heatid="25034" />
                <RESULT resultid="135" eventid="33" swimtime="00:01:09.57" lane="7" heatid="33017" />
                <RESULT resultid="136" eventid="35" swimtime="00:01:19.16" lane="7" heatid="35004" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="28" birthdate="2010-01-01" gender="M" lastname="Piehler" firstname="Junis Arthur" license="408097">
              <RESULTS>
                <RESULT resultid="137" eventid="2" swimtime="00:02:46.29" lane="3" heatid="2007">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:19.89" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="138" eventid="4" swimtime="00:01:24.80" lane="1" heatid="4011" />
                <RESULT resultid="139" eventid="11" swimtime="00:01:23.24" lane="4" heatid="11010" />
                <RESULT resultid="140" eventid="13" swimtime="00:00:31.35" lane="7" heatid="13015" />
                <RESULT resultid="141" eventid="20" swimtime="00:00:39.38" lane="8" heatid="20022" />
                <RESULT resultid="142" eventid="26" swimtime="00:00:38.32" lane="8" heatid="26022" />
                <RESULT resultid="143" eventid="34" swimtime="00:01:11.05" lane="7" heatid="34013" />
                <RESULT resultid="144" eventid="38" swimtime="00:02:51.85" lane="5" heatid="38004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:25.31" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="29" birthdate="2011-01-01" gender="F" lastname="Glatzel" firstname="Lysena" license="418809">
              <RESULTS>
                <RESULT resultid="145" eventid="1" swimtime="00:03:02.43" lane="4" heatid="1004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:28.44" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="146" eventid="3" swimtime="00:01:33.75" lane="8" heatid="3011" />
                <RESULT resultid="147" eventid="10" swimtime="00:01:31.41" lane="5" heatid="10005" />
                <RESULT resultid="148" eventid="14" swimtime="00:03:22.88" lane="5" heatid="14006">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:41.41" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="149" eventid="19" swimtime="00:00:41.17" lane="7" heatid="19025" />
                <RESULT resultid="150" eventid="23" swimtime="00:02:51.26" lane="5" heatid="23006">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:23.98" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="151" eventid="33" swimtime="00:01:20.84" lane="7" heatid="33013" />
                <RESULT resultid="152" eventid="35" swimtime="00:01:34.68" lane="3" heatid="35002" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="30" birthdate="2011-01-01" gender="F" lastname="Forner" firstname="Marleen" license="426142">
              <RESULTS>
                <RESULT resultid="153" eventid="1" swimtime="00:03:01.37" lane="8" heatid="1006">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:25.55" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="154" eventid="5" swimtime="00:00:35.67" lane="7" heatid="5011" />
                <RESULT resultid="155" eventid="10" swimtime="00:01:22.49" lane="5" heatid="10013" />
                <RESULT resultid="156" eventid="12" swimtime="00:00:32.26" lane="1" heatid="12014" />
                <RESULT resultid="157" eventid="19" swimtime="00:00:44.77" lane="7" heatid="19020" />
                <RESULT resultid="158" eventid="23" swimtime="00:02:36.51" lane="3" heatid="23010">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:17.07" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="159" eventid="33" swimtime="00:01:12.66" lane="2" heatid="33014" />
                <RESULT resultid="160" eventid="37" swimtime="00:02:54.87" lane="2" heatid="37007">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:26.30" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="31" birthdate="2012-01-01" gender="M" lastname="Scheinpflug" firstname="Mika" license="445480">
              <RESULTS>
                <RESULT resultid="161" eventid="4" swimtime="00:01:48.82" lane="7" heatid="4005" />
                <RESULT resultid="162" eventid="11" status="DNS" swimtime="00:00:00.00" lane="8" heatid="11004" />
                <RESULT resultid="163" eventid="13" swimtime="00:00:39.71" lane="4" heatid="13006" />
                <RESULT resultid="164" eventid="15" swimtime="00:03:58.73" lane="7" heatid="15003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:58.43" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="165" eventid="20" status="DSQ" swimtime="00:00:50.58" lane="8" heatid="20014" comment="2 Delphinkicks" />
                <RESULT resultid="166" eventid="28" swimtime="00:00:58.75" lane="2" heatid="28008" />
                <RESULT resultid="167" eventid="32" status="DSQ" swimtime="00:01:14.46" lane="8" heatid="32004" comment="Das Brett wurde beim Anschlag nicht vorn umfasst.&#xA;Brustbeinschlag vor dem Ziel." />
                <RESULT resultid="168" eventid="34" swimtime="00:01:36.34" lane="3" heatid="34005" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="32" birthdate="2011-01-01" gender="F" lastname="Schönberg" firstname="Ninett" license="418811">
              <RESULTS>
                <RESULT resultid="169" eventid="3" swimtime="00:01:32.71" lane="5" heatid="3010" />
                <RESULT resultid="170" eventid="5" swimtime="00:00:34.59" lane="6" heatid="5011" />
                <RESULT resultid="171" eventid="10" swimtime="00:01:23.71" lane="7" heatid="10007" />
                <RESULT resultid="172" eventid="12" swimtime="00:00:31.21" lane="6" heatid="12017" />
                <RESULT resultid="173" eventid="19" swimtime="00:00:41.44" lane="1" heatid="19026" />
                <RESULT resultid="174" eventid="25" swimtime="00:00:38.12" lane="6" heatid="25030" />
                <RESULT resultid="175" eventid="33" swimtime="00:01:08.08" lane="6" heatid="33017" />
                <RESULT resultid="176" eventid="35" swimtime="00:01:18.06" lane="2" heatid="35004" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="33" birthdate="2012-01-01" gender="F" lastname="Ballas" firstname="Pauline" license="441075">
              <RESULTS>
                <RESULT resultid="177" eventid="3" swimtime="00:01:39.16" lane="6" heatid="3008" />
                <RESULT resultid="178" eventid="5" swimtime="00:00:42.56" lane="1" heatid="5007" />
                <RESULT resultid="179" eventid="10" swimtime="00:01:29.68" lane="6" heatid="10006" />
                <RESULT resultid="180" eventid="12" swimtime="00:00:35.41" lane="2" heatid="12010" />
                <RESULT resultid="181" eventid="19" swimtime="00:00:45.18" lane="4" heatid="19023" />
                <RESULT resultid="182" eventid="25" swimtime="00:00:42.58" lane="7" heatid="25025" />
                <RESULT resultid="183" eventid="33" swimtime="00:01:16.17" lane="8" heatid="33014" />
                <RESULT resultid="184" eventid="37" swimtime="00:03:09.82" lane="6" heatid="37004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:34.49" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="34" birthdate="2012-01-01" gender="M" lastname="Bodusch" firstname="Tom" license="440974">
              <RESULTS>
                <RESULT resultid="185" eventid="2" swimtime="00:02:49.42" lane="2" heatid="2007">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:15.98" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="186" eventid="6" swimtime="00:00:30.80" lane="7" heatid="6009" />
                <RESULT resultid="187" eventid="11" swimtime="00:01:14.78" lane="4" heatid="11011" />
                <RESULT resultid="188" eventid="13" swimtime="00:00:30.53" lane="2" heatid="13014" />
                <RESULT resultid="189" eventid="22" swimtime="00:00:41.82" lane="4" heatid="22011" />
                <RESULT resultid="190" eventid="26" swimtime="00:00:33.24" lane="2" heatid="26023" />
                <RESULT resultid="191" eventid="32" swimtime="00:00:41.56" lane="4" heatid="32005" />
                <RESULT resultid="192" eventid="34" swimtime="00:01:06.67" lane="6" heatid="34013" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY number="1" gender="X" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="111" eventid="7" swimtime="00:02:15.43" lane="5" heatid="7003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:12.57" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="27" number="1" />
                    <RELAYPOSITION athleteid="28" number="2" />
                    <RELAYPOSITION athleteid="26" number="3" />
                    <RELAYPOSITION athleteid="32" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="2" gender="X" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="112" eventid="7" swimtime="00:02:17.96" lane="6" heatid="7003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:13.79" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="34" number="1" />
                    <RELAYPOSITION athleteid="29" number="2" />
                    <RELAYPOSITION athleteid="25" number="3" />
                    <RELAYPOSITION athleteid="30" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB name="SSV Freiberg" nation="GER" region="12" code="3370">
          <ATHLETES>
            <ATHLETE athleteid="2" birthdate="2013-01-01" gender="F" lastname="Kirchhübel" firstname="Hannah" license="446897">
              <RESULTS>
                <RESULT resultid="7" eventid="1" swimtime="00:03:22.10" lane="2" heatid="1003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:35.40" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="8" eventid="5" swimtime="00:00:39.35" lane="7" heatid="5008" />
                <RESULT resultid="9" eventid="10" swimtime="00:01:32.64" lane="6" heatid="10009" />
                <RESULT resultid="10" eventid="12" swimtime="00:00:36.34" lane="5" heatid="12011" />
                <RESULT resultid="11" eventid="25" swimtime="00:00:39.74" lane="4" heatid="25026" />
                <RESULT resultid="12" eventid="33" swimtime="00:01:25.45" lane="3" heatid="33011" />
                <RESULT resultid="13" eventid="37" swimtime="00:03:18.28" lane="3" heatid="37004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:37.40" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="3" birthdate="2012-01-01" gender="F" lastname="Lampke" firstname="Ingrid" license="433827">
              <RESULTS>
                <RESULT resultid="14" eventid="1" swimtime="00:03:07.80" lane="1" heatid="1004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:30.14" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="15" eventid="5" swimtime="00:00:35.79" lane="6" heatid="5009" />
                <RESULT resultid="16" eventid="10" swimtime="00:01:28.05" lane="2" heatid="10011" />
                <RESULT resultid="17" eventid="12" swimtime="00:00:31.95" lane="6" heatid="12014" />
                <RESULT resultid="18" eventid="23" swimtime="00:02:49.27" lane="8" heatid="23009">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:23.03" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="19" eventid="25" swimtime="00:00:40.30" lane="4" heatid="25027" />
                <RESULT resultid="20" eventid="33" swimtime="00:01:15.14" lane="1" heatid="33013" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="4" birthdate="2011-01-01" gender="F" lastname="Emmrich" firstname="Leonie" license="421842">
              <RESULTS>
                <RESULT resultid="21" eventid="23" swimtime="00:02:44.08" lane="5" heatid="23007">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:17.49" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="22" eventid="25" swimtime="00:00:38.94" lane="1" heatid="25032" />
                <RESULT resultid="23" eventid="33" swimtime="00:01:13.81" lane="1" heatid="33015" />
                <RESULT resultid="24" eventid="37" swimtime="00:03:11.80" lane="8" heatid="37005">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:34.31" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="SSV Hoyerswerda" nation="GER" region="12" code="3374">
          <ATHLETES>
            <ATHLETE athleteid="976" birthdate="2014-01-01" gender="M" lastname="Steyreiff" firstname="Anton" license="465606">
              <RESULTS>
                <RESULT resultid="4532" eventid="18" swimtime="00:01:03.20" lane="4" heatid="18009" />
                <RESULT resultid="4533" eventid="20" swimtime="00:00:59.96" lane="7" heatid="20008" />
                <RESULT resultid="4534" eventid="28" swimtime="00:01:06.73" lane="3" heatid="28001" />
                <RESULT resultid="4535" eventid="30" swimtime="00:00:51.36" lane="3" heatid="30003" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="977" birthdate="2009-01-01" gender="M" lastname="Szczepanski" firstname="Benjamin" license="402425">
              <RESULTS>
                <RESULT resultid="4536" eventid="4" swimtime="00:01:41.70" lane="1" heatid="4007" />
                <RESULT resultid="4537" eventid="13" swimtime="00:00:37.06" lane="5" heatid="13004" />
                <RESULT resultid="4538" eventid="20" swimtime="00:00:44.87" lane="5" heatid="20015" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="978" birthdate="2010-01-01" gender="M" lastname="Puls" firstname="Dennis" license="411461">
              <RESULTS>
                <RESULT resultid="4539" eventid="6" swimtime="00:00:52.93" lane="7" heatid="6001" />
                <RESULT resultid="4540" eventid="11" swimtime="00:01:36.97" lane="7" heatid="11005" />
                <RESULT resultid="4541" eventid="13" swimtime="00:00:36.19" lane="8" heatid="13008" />
                <RESULT resultid="4542" eventid="24" swimtime="00:03:01.65" lane="1" heatid="24002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:24.39" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="4543" eventid="26" swimtime="00:00:43.23" lane="1" heatid="26017" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="979" birthdate="2011-01-01" gender="F" lastname="Schädrich" firstname="Emma" license="426979">
              <RESULTS>
                <RESULT resultid="4544" eventid="1" swimtime="00:03:27.26" lane="7" heatid="1002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:36.46" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="4545" eventid="3" swimtime="00:01:40.90" lane="7" heatid="3007" />
                <RESULT resultid="4546" eventid="12" swimtime="00:00:35.54" lane="2" heatid="12011" />
                <RESULT resultid="4547" eventid="14" swimtime="00:03:39.34" lane="7" heatid="14004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:44.16" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="4548" eventid="19" swimtime="00:00:43.46" lane="7" heatid="19024" />
                <RESULT resultid="4549" eventid="23" swimtime="00:03:03.96" lane="6" heatid="23002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:30.69" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="4550" eventid="25" swimtime="00:00:42.09" lane="3" heatid="25024" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="980" birthdate="2010-01-01" gender="M" lastname="Korch" firstname="Fabian" license="422439">
              <RESULTS>
                <RESULT resultid="4551" eventid="4" swimtime="00:01:37.33" lane="3" heatid="4005" />
                <RESULT resultid="4552" eventid="13" swimtime="00:00:35.41" lane="7" heatid="13008" />
                <RESULT resultid="4553" eventid="15" status="DSQ" swimtime="00:03:37.67" lane="5" heatid="15001" comment="Anschlag an der 3. Wende mit einer Hand.">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:44.96" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="4554" eventid="20" swimtime="00:00:42.11" lane="6" heatid="20018" />
                <RESULT resultid="4555" eventid="26" swimtime="00:00:45.67" lane="2" heatid="26015" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="981" birthdate="2011-01-01" gender="F" lastname="Szczepanski" firstname="Helena" license="425743">
              <RESULTS>
                <RESULT resultid="4556" eventid="5" swimtime="00:00:49.78" lane="3" heatid="5004" />
                <RESULT resultid="4557" eventid="10" swimtime="00:01:41.35" lane="5" heatid="10003" />
                <RESULT resultid="4558" eventid="12" swimtime="00:00:41.05" lane="2" heatid="12004" />
                <RESULT resultid="4559" eventid="19" swimtime="00:00:55.83" lane="1" heatid="19012" />
                <RESULT resultid="4560" eventid="25" swimtime="00:00:45.10" lane="5" heatid="25021" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="982" birthdate="2012-01-01" gender="F" lastname="Grosa" firstname="Helene" license="460071">
              <RESULTS>
                <RESULT resultid="4561" eventid="19" swimtime="00:00:54.86" lane="5" heatid="19013" />
                <RESULT resultid="4562" eventid="25" swimtime="00:00:54.63" lane="1" heatid="25012" />
                <RESULT resultid="4563" eventid="27" swimtime="00:01:07.48" lane="8" heatid="27002" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="983" birthdate="2010-01-01" gender="M" lastname="Grosa" firstname="Johann" license="425731">
              <RESULTS>
                <RESULT resultid="4564" eventid="20" status="DSQ" swimtime="00:00:44.68" lane="4" heatid="20016" comment="Start vor dem Startsignal." />
                <RESULT resultid="4565" eventid="24" swimtime="00:03:01.08" lane="3" heatid="24001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:26.26" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="4566" eventid="26" swimtime="00:00:47.30" lane="5" heatid="26011" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="984" birthdate="2010-01-01" gender="M" lastname="Schneider" firstname="Johannes" license="416453">
              <RESULTS>
                <RESULT resultid="4567" eventid="4" swimtime="00:01:45.47" lane="3" heatid="4002" />
                <RESULT resultid="4568" eventid="6" status="DSQ" swimtime="00:00:54.87" lane="8" heatid="6004" comment="Schwimmer beendete die Schwimmstrecke mit Brustschwimmen." />
                <RESULT resultid="4569" eventid="11" swimtime="00:01:46.84" lane="6" heatid="11004" />
                <RESULT resultid="4570" eventid="13" swimtime="00:00:37.35" lane="6" heatid="13005" />
                <RESULT resultid="4571" eventid="20" swimtime="00:00:46.06" lane="4" heatid="20013" />
                <RESULT resultid="4572" eventid="26" swimtime="00:00:43.64" lane="2" heatid="26014" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="985" birthdate="2007-01-01" gender="M" lastname="Püschel" firstname="Jonas" license="376888">
              <RESULTS>
                <RESULT resultid="4573" eventid="2" swimtime="00:02:40.25" lane="8" heatid="2007">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:10.42" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="4574" eventid="6" swimtime="00:00:28.44" lane="2" heatid="6011" />
                <RESULT resultid="4575" eventid="11" swimtime="00:01:11.69" lane="1" heatid="11012" />
                <RESULT resultid="4576" eventid="13" swimtime="00:00:27.06" lane="7" heatid="13018" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="986" birthdate="2008-01-01" gender="F" lastname="Senf" firstname="Leonie" license="388279">
              <RESULTS>
                <RESULT resultid="4577" eventid="1" swimtime="00:02:46.07" lane="2" heatid="1007">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:18.85" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="4578" eventid="5" swimtime="00:00:31.45" lane="4" heatid="5013" />
                <RESULT resultid="4579" eventid="10" swimtime="00:01:16.89" lane="8" heatid="10016" />
                <RESULT resultid="4580" eventid="12" swimtime="00:00:30.25" lane="2" heatid="12018" />
                <RESULT resultid="4581" eventid="19" swimtime="00:00:37.54" lane="4" heatid="19026" />
                <RESULT resultid="4582" eventid="23" swimtime="00:02:28.65" lane="3" heatid="23011">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:09.63" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="4583" eventid="25" swimtime="00:00:34.96" lane="7" heatid="25034" />
                <RESULT resultid="4584" eventid="33" swimtime="00:01:05.74" lane="6" heatid="33018" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="987" birthdate="2015-01-01" gender="F" lastname="Modsching" firstname="Lucy Jolene" license="465612">
              <RESULTS>
                <RESULT resultid="4585" eventid="19" swimtime="00:00:54.61" lane="2" heatid="19010" />
                <RESULT resultid="4586" eventid="21" swimtime="00:01:07.10" lane="4" heatid="21001" />
                <RESULT resultid="4587" eventid="25" swimtime="00:01:05.14" lane="4" heatid="25005" />
                <RESULT resultid="4588" eventid="27" swimtime="00:01:06.50" lane="1" heatid="27009" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="988" birthdate="2010-01-01" gender="M" lastname="Seeger" firstname="Quin" license="432231">
              <RESULTS>
                <RESULT resultid="4589" eventid="2" swimtime="00:03:09.77" lane="2" heatid="2003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:31.99" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="4590" eventid="6" swimtime="00:00:36.64" lane="7" heatid="6007" />
                <RESULT resultid="4591" eventid="11" swimtime="00:01:36.48" lane="8" heatid="11003" />
                <RESULT resultid="4592" eventid="13" swimtime="00:00:30.66" lane="6" heatid="13014" />
                <RESULT resultid="4593" eventid="20" swimtime="00:00:42.34" lane="8" heatid="20019" />
                <RESULT resultid="4594" eventid="24" swimtime="00:02:43.30" lane="6" heatid="24003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:17.82" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="4595" eventid="26" status="DSQ" swimtime="00:00:39.73" lane="7" heatid="26020" comment="Start vor dem Startsignal." />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="989" birthdate="2009-01-01" gender="M" lastname="Janze" firstname="Roque" license="399802">
              <RESULTS>
                <RESULT resultid="4596" eventid="4" swimtime="00:01:31.71" lane="7" heatid="4008" />
                <RESULT resultid="4597" eventid="11" swimtime="00:01:19.20" lane="3" heatid="11009" />
                <RESULT resultid="4598" eventid="13" swimtime="00:00:33.45" lane="6" heatid="13012" />
                <RESULT resultid="4599" eventid="15" swimtime="00:03:29.78" lane="4" heatid="15004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:43.43" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="4600" eventid="20" swimtime="00:00:40.08" lane="6" heatid="20019" />
                <RESULT resultid="4601" eventid="24" swimtime="00:02:45.89" lane="2" heatid="24002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:19.51" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="4602" eventid="26" swimtime="00:00:36.77" lane="3" heatid="26022" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="990" birthdate="2011-01-01" gender="M" lastname="Dzikowski" firstname="Theo" license="460074">
              <RESULTS>
                <RESULT resultid="4603" eventid="6" swimtime="00:00:41.92" lane="7" heatid="6004" />
                <RESULT resultid="4604" eventid="11" swimtime="00:01:38.52" lane="6" heatid="11003" />
                <RESULT resultid="4605" eventid="13" swimtime="00:00:34.59" lane="1" heatid="13009" />
                <RESULT resultid="4606" eventid="24" swimtime="00:02:55.07" lane="6" heatid="24001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:24.14" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="4607" eventid="26" swimtime="00:00:44.36" lane="8" heatid="26016" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="991" birthdate="2010-01-01" gender="M" lastname="Hoffmann" firstname="Valentin" license="416450">
              <RESULTS>
                <RESULT resultid="4608" eventid="6" swimtime="00:00:43.26" lane="5" heatid="6003" />
                <RESULT resultid="4609" eventid="11" swimtime="00:01:42.70" lane="3" heatid="11005" />
                <RESULT resultid="4610" eventid="13" swimtime="00:00:36.45" lane="8" heatid="13009" />
                <RESULT resultid="4611" eventid="24" swimtime="00:03:10.32" lane="8" heatid="24002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:27.63" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="4612" eventid="26" swimtime="00:00:45.49" lane="6" heatid="26015" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY number="1" gender="X" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="4530" eventid="16" swimtime="00:02:20.68" lane="4" heatid="16001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:22.32" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="989" number="1" />
                    <RELAYPOSITION athleteid="977" number="2" />
                    <RELAYPOSITION athleteid="985" number="3" />
                    <RELAYPOSITION athleteid="986" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" gender="X" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="4531" eventid="7" swimtime="00:02:37.55" lane="5" heatid="7002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:25.08" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="978" number="1" />
                    <RELAYPOSITION athleteid="980" number="2" />
                    <RELAYPOSITION athleteid="988" number="3" />
                    <RELAYPOSITION athleteid="979" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB name="SSV Leutzsch" nation="GER" region="12" code="3378">
          <ATHLETES>
            <ATHLETE athleteid="155" birthdate="2012-01-01" gender="M" lastname="Kotliarov" firstname="Albert" license="475776">
              <RESULTS>
                <RESULT resultid="816" eventid="6" swimtime="00:00:48.95" lane="8" heatid="6001" />
                <RESULT resultid="815" eventid="11" status="DSQ" swimtime="00:01:41.34" lane="3" heatid="11001" comment="Hat sich bei der Wende nicht in Rückenlage abgestoßen." />
                <RESULT resultid="814" eventid="13" swimtime="00:00:37.75" lane="4" heatid="13004" />
                <RESULT resultid="813" eventid="18" swimtime="00:01:01.72" lane="7" heatid="18009" />
                <RESULT resultid="812" eventid="24" swimtime="00:03:10.09" lane="4" heatid="24001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:29.03" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="811" eventid="34" status="DNS" swimtime="00:00:00.00" lane="6" heatid="34005" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="156" birthdate="2012-01-01" gender="M" lastname="Khrushch" firstname="Yakiv" license="429613">
              <RESULTS>
                <RESULT resultid="824" eventid="2" swimtime="00:02:56.39" lane="2" heatid="2006">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:24.03" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="823" eventid="4" swimtime="00:01:36.99" lane="5" heatid="4007" />
                <RESULT resultid="822" eventid="11" swimtime="00:01:21.50" lane="8" heatid="11010" />
                <RESULT resultid="821" eventid="15" swimtime="00:03:25.82" lane="8" heatid="15005">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:40.27" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="820" eventid="20" swimtime="00:00:44.34" lane="2" heatid="20017" />
                <RESULT resultid="819" eventid="26" swimtime="00:00:39.00" lane="5" heatid="26020" />
                <RESULT resultid="818" eventid="34" swimtime="00:01:12.65" lane="8" heatid="34012" />
                <RESULT resultid="817" eventid="38" swimtime="00:02:54.16" lane="3" heatid="38004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:27.42" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="157" birthdate="2013-01-01" gender="M" lastname="Plewa" firstname="Valentin" license="441003">
              <RESULTS>
                <RESULT resultid="831" eventid="2" swimtime="00:03:14.67" lane="5" heatid="2004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:33.27" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="830" eventid="6" swimtime="00:00:36.79" lane="1" heatid="6007" />
                <RESULT resultid="829" eventid="13" swimtime="00:00:36.84" lane="3" heatid="13006" />
                <RESULT resultid="828" eventid="20" status="DNS" swimtime="00:00:00.00" lane="6" heatid="20013" />
                <RESULT resultid="827" eventid="24" status="DNS" swimtime="00:00:00.00" lane="8" heatid="24004" />
                <RESULT resultid="826" eventid="28" status="DNS" swimtime="00:00:00.00" lane="8" heatid="28008" />
                <RESULT resultid="825" eventid="34" status="DNS" swimtime="00:00:00.00" lane="6" heatid="34008" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="158" birthdate="2015-01-01" gender="M" lastname="Albert" firstname="Theo" license="466653">
              <RESULTS>
                <RESULT resultid="834" eventid="18" swimtime="00:01:17.88" lane="2" heatid="18003" />
                <RESULT resultid="833" eventid="26" swimtime="00:01:04.07" lane="7" heatid="26003" />
                <RESULT resultid="832" eventid="30" swimtime="00:01:06.62" lane="6" heatid="30001" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="159" birthdate="2014-01-01" gender="F" lastname="Richter" firstname="Stella" license="466191">
              <RESULTS>
                <RESULT resultid="839" eventid="17" swimtime="00:01:16.67" lane="4" heatid="17004" />
                <RESULT resultid="838" eventid="21" swimtime="00:01:19.47" lane="5" heatid="21002" />
                <RESULT resultid="837" eventid="25" swimtime="00:01:04.96" lane="3" heatid="25002" />
                <RESULT resultid="836" eventid="29" swimtime="00:00:58.01" lane="1" heatid="29003" />
                <RESULT resultid="835" eventid="31" swimtime="00:01:27.52" lane="3" heatid="31001" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="160" birthdate="2013-01-01" gender="F" lastname="Riemer" firstname="Sonja" license="461030">
              <RESULTS>
                <RESULT resultid="846" eventid="1" swimtime="00:03:36.85" lane="1" heatid="1002" />
                <RESULT resultid="845" eventid="5" swimtime="00:00:41.29" lane="6" heatid="5005" />
                <RESULT resultid="844" eventid="10" swimtime="00:01:41.96" lane="8" heatid="10005" />
                <RESULT resultid="843" eventid="12" swimtime="00:00:38.76" lane="8" heatid="12004" />
                <RESULT resultid="842" eventid="17" swimtime="00:01:06.53" lane="4" heatid="17003" />
                <RESULT resultid="841" eventid="21" swimtime="00:00:57.44" lane="6" heatid="21011" />
                <RESULT resultid="840" eventid="23" swimtime="00:03:10.45" lane="5" heatid="23002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:32.68" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="161" birthdate="2013-01-01" gender="M" lastname="Kolonko" firstname="Rèmy" license="446750">
              <RESULTS>
                <RESULT resultid="853" eventid="4" swimtime="00:01:40.74" lane="6" heatid="4007" />
                <RESULT resultid="852" eventid="13" swimtime="00:00:36.18" lane="8" heatid="13006" />
                <RESULT resultid="851" eventid="15" swimtime="00:03:43.21" lane="3" heatid="15003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:50.74" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="850" eventid="20" swimtime="00:00:44.39" lane="5" heatid="20016" />
                <RESULT resultid="849" eventid="28" swimtime="00:00:55.00" lane="6" heatid="28008" />
                <RESULT resultid="848" eventid="32" swimtime="00:01:00.53" lane="3" heatid="32004" />
                <RESULT resultid="847" eventid="34" swimtime="00:01:25.79" lane="1" heatid="34006" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="162" birthdate="2012-01-01" gender="M" lastname="Fabricius" firstname="Paul" license="443229">
              <RESULTS>
                <RESULT resultid="860" eventid="4" swimtime="00:01:59.10" lane="6" heatid="4002" />
                <RESULT resultid="859" eventid="11" swimtime="00:01:39.51" lane="5" heatid="11004" />
                <RESULT resultid="858" eventid="13" swimtime="00:00:40.22" lane="8" heatid="13005" />
                <RESULT resultid="857" eventid="18" swimtime="00:01:07.24" lane="2" heatid="18005" />
                <RESULT resultid="856" eventid="24" swimtime="00:03:09.48" lane="2" heatid="24003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:33.68" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="855" eventid="34" swimtime="00:01:28.54" lane="4" heatid="34005" />
                <RESULT resultid="854" eventid="38" swimtime="00:03:26.31" lane="7" heatid="38001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:42.21" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="163" birthdate="2015-01-01" gender="M" lastname="Laut" firstname="Oliver Alexander" license="463402">
              <RESULTS>
                <RESULT resultid="864" eventid="18" swimtime="00:01:13.19" lane="7" heatid="18005" />
                <RESULT resultid="863" eventid="20" swimtime="00:01:06.20" lane="3" heatid="20004" />
                <RESULT resultid="862" eventid="28" swimtime="00:01:05.84" lane="5" heatid="28005" />
                <RESULT resultid="861" eventid="30" swimtime="00:01:00.48" lane="2" heatid="30002" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="164" birthdate="2015-01-01" gender="F" lastname="Schüler" firstname="Mila" license="463401">
              <RESULTS>
                <RESULT resultid="868" eventid="17" swimtime="00:01:16.03" lane="6" heatid="17003" />
                <RESULT resultid="867" eventid="21" swimtime="00:01:18.17" lane="1" heatid="21003" />
                <RESULT resultid="866" eventid="25" swimtime="00:01:05.50" lane="6" heatid="25004" />
                <RESULT resultid="865" eventid="29" swimtime="00:01:06.73" lane="4" heatid="29001" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="165" birthdate="2010-01-01" gender="M" lastname="Leonhardt" firstname="Mika" license="405569">
              <RESULTS>
                <RESULT resultid="875" eventid="2" swimtime="00:02:38.83" lane="8" heatid="2008">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:14.14" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="874" eventid="6" swimtime="00:00:30.76" lane="8" heatid="6011" />
                <RESULT resultid="873" eventid="9" swimtime="00:02:39.00" lane="4" heatid="9001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:13.65" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="872" eventid="13" swimtime="00:00:29.39" lane="1" heatid="13016" />
                <RESULT resultid="871" eventid="20" swimtime="00:00:38.99" lane="2" heatid="20018" />
                <RESULT resultid="870" eventid="24" swimtime="00:02:21.91" lane="3" heatid="24008">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:10.05" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="869" eventid="36" swimtime="00:01:11.37" lane="3" heatid="36003" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="166" birthdate="2015-01-01" gender="F" lastname="Markov" firstname="Mathilda" license="463355">
              <RESULTS>
                <RESULT resultid="879" eventid="17" swimtime="00:01:03.52" lane="1" heatid="17013" />
                <RESULT resultid="878" eventid="21" swimtime="00:00:58.65" lane="8" heatid="21009" />
                <RESULT resultid="877" eventid="25" swimtime="00:00:53.50" lane="6" heatid="25014" />
                <RESULT resultid="876" eventid="29" swimtime="00:00:50.69" lane="5" heatid="29006" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="167" birthdate="2014-01-01" gender="M" lastname="Jung" firstname="Mateo" license="446744">
              <RESULTS>
                <RESULT resultid="884" eventid="18" swimtime="00:00:53.93" lane="4" heatid="18011" />
                <RESULT resultid="883" eventid="22" swimtime="00:00:48.53" lane="3" heatid="22011" />
                <RESULT resultid="882" eventid="26" swimtime="00:00:46.66" lane="3" heatid="26016" />
                <RESULT resultid="881" eventid="30" swimtime="00:00:39.82" lane="3" heatid="30008" />
                <RESULT resultid="880" eventid="32" swimtime="00:00:58.93" lane="1" heatid="32005" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="168" birthdate="2013-01-01" gender="F" lastname="Frank" firstname="Martha Leni" license="441008">
              <RESULTS>
                <RESULT resultid="891" eventid="5" swimtime="00:00:39.91" lane="3" heatid="5006" />
                <RESULT resultid="890" eventid="10" swimtime="00:01:33.29" lane="5" heatid="10008" />
                <RESULT resultid="889" eventid="12" swimtime="00:00:36.79" lane="8" heatid="12008" />
                <RESULT resultid="888" eventid="17" swimtime="00:00:53.32" lane="4" heatid="17013" />
                <RESULT resultid="887" eventid="21" swimtime="00:00:54.42" lane="5" heatid="21013" />
                <RESULT resultid="886" eventid="25" swimtime="00:00:43.35" lane="8" heatid="25026" />
                <RESULT resultid="885" eventid="31" swimtime="00:00:56.69" lane="1" heatid="31007" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="169" birthdate="2013-01-01" gender="F" lastname="Petzold" firstname="Malin" license="445609">
              <RESULTS>
                <RESULT resultid="898" eventid="3" swimtime="00:01:44.93" lane="7" heatid="3006" />
                <RESULT resultid="897" eventid="12" swimtime="00:00:39.12" lane="1" heatid="12008" />
                <RESULT resultid="896" eventid="14" swimtime="00:03:50.74" lane="1" heatid="14005">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:51.80" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="895" eventid="19" status="WDR" swimtime="00:00:00.00" lane="2" heatid="19022" />
                <RESULT resultid="894" eventid="27" status="WDR" swimtime="00:00:00.00" lane="1" heatid="27012" />
                <RESULT resultid="893" eventid="33" status="WDR" swimtime="00:00:00.00" lane="8" heatid="33011" />
                <RESULT resultid="892" eventid="37" status="WDR" swimtime="00:00:00.00" lane="4" heatid="37002" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="170" birthdate="2015-01-01" gender="F" lastname="Herold" firstname="Lotta" license="466193">
              <RESULTS>
                <RESULT resultid="902" eventid="19" swimtime="00:01:03.31" lane="2" heatid="19001" />
                <RESULT resultid="901" eventid="25" swimtime="00:01:02.98" lane="4" heatid="25004" />
                <RESULT resultid="900" eventid="27" swimtime="00:01:13.45" lane="8" heatid="27007" />
                <RESULT resultid="899" eventid="29" swimtime="00:01:15.27" lane="3" heatid="29001" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="171" birthdate="2015-01-01" gender="F" lastname="Kaltenbach" firstname="Livia" license="463353">
              <RESULTS>
                <RESULT resultid="906" eventid="19" swimtime="00:01:01.31" lane="3" heatid="19007" />
                <RESULT resultid="905" eventid="25" swimtime="00:01:02.17" lane="7" heatid="25008" />
                <RESULT resultid="904" eventid="27" swimtime="00:01:13.48" lane="2" heatid="27003" />
                <RESULT resultid="903" eventid="29" swimtime="00:00:54.20" lane="7" heatid="29005" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="172" birthdate="2014-01-01" gender="F" lastname="Schuster" firstname="Lina-Collien" license="466282">
              <RESULTS>
                <RESULT resultid="911" eventid="17" swimtime="00:01:01.68" lane="3" heatid="17010" />
                <RESULT resultid="910" eventid="25" swimtime="00:00:53.70" lane="2" heatid="25011" />
                <RESULT resultid="909" eventid="29" swimtime="00:00:47.83" lane="6" heatid="29006" />
                <RESULT resultid="908" eventid="31" swimtime="00:01:05.08" lane="4" heatid="31003" />
                <RESULT resultid="907" eventid="33" swimtime="00:01:46.26" lane="5" heatid="33001" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="173" birthdate="2012-01-01" gender="M" lastname="Seifert" firstname="Leo Arend" license="444237">
              <RESULTS>
                <RESULT resultid="918" eventid="6" swimtime="00:00:39.71" lane="4" heatid="6006" />
                <RESULT resultid="917" eventid="11" swimtime="00:01:34.29" lane="8" heatid="11007" />
                <RESULT resultid="916" eventid="13" swimtime="00:00:33.88" lane="4" heatid="13010" />
                <RESULT resultid="915" eventid="24" swimtime="00:02:52.40" lane="5" heatid="24005">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:23.72" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="914" eventid="26" swimtime="00:00:42.48" lane="4" heatid="26015" />
                <RESULT resultid="913" eventid="34" swimtime="00:01:16.70" lane="8" heatid="34010" />
                <RESULT resultid="912" eventid="38" swimtime="00:03:18.03" lane="6" heatid="38002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:36.67" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="174" birthdate="2014-01-01" gender="F" lastname="Miemczyk" firstname="Lamiah Soey" license="446742">
              <RESULTS>
                <RESULT resultid="923" eventid="19" swimtime="00:00:54.36" lane="1" heatid="19013" />
                <RESULT resultid="922" eventid="21" swimtime="00:01:02.58" lane="8" heatid="21010" />
                <RESULT resultid="921" eventid="27" swimtime="00:01:03.45" lane="5" heatid="27006" />
                <RESULT resultid="920" eventid="29" swimtime="00:00:44.23" lane="3" heatid="29010" />
                <RESULT resultid="919" eventid="31" swimtime="00:01:02.63" lane="6" heatid="31004" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="175" birthdate="2014-01-01" gender="M" lastname="Keil" firstname="Konrad" license="451443">
              <RESULTS>
                <RESULT resultid="927" eventid="20" swimtime="00:00:56.94" lane="4" heatid="20007" />
                <RESULT resultid="926" eventid="26" swimtime="00:00:59.87" lane="6" heatid="26005" />
                <RESULT resultid="925" eventid="28" swimtime="00:01:05.21" lane="1" heatid="28005" />
                <RESULT resultid="924" eventid="30" swimtime="00:00:51.09" lane="1" heatid="30004" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="176" birthdate="2015-01-01" gender="M" lastname="Haupt" firstname="Konrad Arthur" license="463404">
              <RESULTS>
                <RESULT resultid="931" eventid="20" swimtime="00:01:07.83" lane="2" heatid="20001" />
                <RESULT resultid="930" eventid="26" swimtime="00:01:04.58" lane="8" heatid="26003" />
                <RESULT resultid="929" eventid="28" swimtime="00:01:26.12" lane="1" heatid="28002" />
                <RESULT resultid="928" eventid="30" swimtime="00:01:05.77" lane="7" heatid="30001" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="177" birthdate="2014-01-01" gender="F" lastname="Soto Drewniak" firstname="Klara Filippa" license="466186">
              <RESULTS>
                <RESULT resultid="936" eventid="19" swimtime="00:00:55.80" lane="4" heatid="19012" />
                <RESULT resultid="935" eventid="25" swimtime="00:00:49.85" lane="5" heatid="25015" />
                <RESULT resultid="934" eventid="27" swimtime="00:01:00.24" lane="8" heatid="27011" />
                <RESULT resultid="933" eventid="29" swimtime="00:00:51.61" lane="8" heatid="29007" />
                <RESULT resultid="932" eventid="31" swimtime="00:01:10.23" lane="5" heatid="31003" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="178" birthdate="2015-01-01" gender="M" lastname="Fischer" firstname="Johan" license="473958">
              <RESULTS>
                <RESULT resultid="940" eventid="18" swimtime="00:01:21.25" lane="1" heatid="18003" />
                <RESULT resultid="939" eventid="22" swimtime="00:01:07.47" lane="8" heatid="22002" />
                <RESULT resultid="938" eventid="26" swimtime="00:00:57.11" lane="2" heatid="26002" />
                <RESULT resultid="937" eventid="30" swimtime="00:00:58.96" lane="8" heatid="30001" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="179" birthdate="2013-01-01" gender="M" lastname="Müller" firstname="Jasper" license="441004">
              <RESULTS>
                <RESULT resultid="946" eventid="6" swimtime="00:00:38.75" lane="5" heatid="6004" />
                <RESULT resultid="945" eventid="11" swimtime="00:01:27.81" lane="7" heatid="11009" />
                <RESULT resultid="944" eventid="13" swimtime="00:00:35.39" lane="2" heatid="13011" />
                <RESULT resultid="943" eventid="26" swimtime="00:00:39.27" lane="8" heatid="26021" />
                <RESULT resultid="942" eventid="34" swimtime="00:01:20.52" lane="8" heatid="34009" />
                <RESULT resultid="941" eventid="38" swimtime="00:03:04.81" lane="8" heatid="38004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:32.19" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="180" birthdate="2013-01-01" gender="F" lastname="Ringel" firstname="Ida Emilia" license="446748">
              <RESULTS>
                <RESULT resultid="953" eventid="5" swimtime="00:00:57.40" lane="5" heatid="5001" />
                <RESULT resultid="952" eventid="10" swimtime="00:01:54.08" lane="2" heatid="10002" />
                <RESULT resultid="951" eventid="12" swimtime="00:00:56.63" lane="1" heatid="12002" />
                <RESULT resultid="950" eventid="17" swimtime="00:01:09.52" lane="8" heatid="17007" />
                <RESULT resultid="949" eventid="21" swimtime="00:01:07.75" lane="5" heatid="21007" />
                <RESULT resultid="948" eventid="25" swimtime="00:00:54.37" lane="8" heatid="25013" />
                <RESULT resultid="947" eventid="31" swimtime="00:01:10.03" lane="2" heatid="31004" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="181" birthdate="2012-01-01" gender="F" lastname="Haupt" firstname="Helena Sophie" license="443234">
              <RESULTS>
                <RESULT resultid="961" eventid="3" swimtime="00:01:38.16" lane="1" heatid="3007" />
                <RESULT resultid="960" eventid="5" swimtime="00:00:37.59" lane="2" heatid="5009" />
                <RESULT resultid="959" eventid="10" swimtime="00:01:29.11" lane="6" heatid="10011" />
                <RESULT resultid="958" eventid="12" swimtime="00:00:32.51" lane="6" heatid="12015" />
                <RESULT resultid="957" eventid="17" swimtime="00:00:48.16" lane="2" heatid="17016" />
                <RESULT resultid="956" eventid="25" swimtime="00:00:38.59" lane="3" heatid="25032" />
                <RESULT resultid="955" eventid="33" swimtime="00:01:13.50" lane="6" heatid="33015" />
                <RESULT resultid="954" eventid="37" swimtime="00:03:14.16" lane="2" heatid="37004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:37.55" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="182" birthdate="2014-01-01" gender="F" lastname="Leonhardt" firstname="Hanna" license="446794">
              <RESULTS>
                <RESULT resultid="966" eventid="17" swimtime="00:00:55.02" lane="8" heatid="17016" />
                <RESULT resultid="965" eventid="25" swimtime="00:00:41.69" lane="2" heatid="25028" />
                <RESULT resultid="964" eventid="29" swimtime="00:00:36.12" lane="4" heatid="29013" />
                <RESULT resultid="963" eventid="31" swimtime="00:00:53.19" lane="4" heatid="31006" />
                <RESULT resultid="962" eventid="33" swimtime="00:01:23.89" lane="5" heatid="33011" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="183" birthdate="2015-01-01" gender="M" lastname="Schlott" firstname="Gustav" license="463334">
              <RESULTS>
                <RESULT resultid="970" eventid="18" swimtime="00:01:16.08" lane="8" heatid="18006" />
                <RESULT resultid="969" eventid="22" swimtime="00:01:09.95" lane="3" heatid="22004" />
                <RESULT resultid="968" eventid="26" swimtime="00:00:52.64" lane="3" heatid="26006" />
                <RESULT resultid="967" eventid="30" swimtime="00:00:49.05" lane="2" heatid="30004" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="184" birthdate="2011-01-01" gender="F" lastname="Reyher" firstname="Frida Emily" license="423155">
              <RESULTS>
                <RESULT resultid="978" eventid="1" swimtime="00:02:56.87" lane="3" heatid="1006">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:23.73" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="977" eventid="5" swimtime="00:00:38.70" lane="8" heatid="5009" />
                <RESULT resultid="976" eventid="10" swimtime="00:01:21.59" lane="7" heatid="10015" />
                <RESULT resultid="975" eventid="12" swimtime="00:00:33.45" lane="8" heatid="12015" />
                <RESULT resultid="974" eventid="23" swimtime="00:02:32.48" lane="8" heatid="23011">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:14.30" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="973" eventid="25" swimtime="00:00:36.17" lane="6" heatid="25033" />
                <RESULT resultid="972" eventid="33" swimtime="00:01:12.52" lane="1" heatid="33016" />
                <RESULT resultid="971" eventid="37" swimtime="00:02:50.99" lane="6" heatid="37007">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:25.28" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="185" birthdate="2014-01-01" gender="M" lastname="Ronneberger" firstname="Djamel" license="451441">
              <RESULTS>
                <RESULT resultid="983" eventid="18" swimtime="00:01:00.79" lane="4" heatid="18007" />
                <RESULT resultid="982" eventid="20" status="DSQ" swimtime="00:01:01.62" lane="2" heatid="20004" comment="mehrere Kraulbeinschläge nach dem Start." />
                <RESULT resultid="981" eventid="26" swimtime="00:00:54.33" lane="5" heatid="26005" />
                <RESULT resultid="980" eventid="28" swimtime="00:01:11.29" lane="3" heatid="28003" />
                <RESULT resultid="979" eventid="30" swimtime="00:00:58.53" lane="3" heatid="30001" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="186" birthdate="2014-01-01" gender="M" lastname="Mönch" firstname="Darwin" license="458348">
              <RESULTS>
                <RESULT resultid="987" eventid="20" swimtime="00:01:02.48" lane="4" heatid="20003" />
                <RESULT resultid="986" eventid="26" swimtime="00:01:02.40" lane="3" heatid="26003" />
                <RESULT resultid="985" eventid="28" swimtime="00:01:12.02" lane="5" heatid="28003" />
                <RESULT resultid="984" eventid="30" swimtime="00:01:07.24" lane="5" heatid="30001" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="187" birthdate="2012-01-01" gender="M" lastname="Aprodu" firstname="Daniil" license="438637">
              <RESULTS>
                <RESULT resultid="995" eventid="2" swimtime="00:03:27.39" lane="4" heatid="2003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:37.27" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="994" eventid="6" swimtime="00:00:42.87" lane="4" heatid="6003" />
                <RESULT resultid="993" eventid="11" swimtime="00:01:36.43" lane="2" heatid="11006" />
                <RESULT resultid="992" eventid="13" swimtime="00:00:36.51" lane="3" heatid="13008" />
                <RESULT resultid="991" eventid="18" swimtime="00:01:01.09" lane="1" heatid="18011" />
                <RESULT resultid="990" eventid="24" swimtime="00:03:01.57" lane="6" heatid="24004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:27.58" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="989" eventid="34" swimtime="00:01:23.46" lane="8" heatid="34008" />
                <RESULT resultid="988" eventid="38" swimtime="00:03:18.55" lane="7" heatid="38002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:38.75" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="188" birthdate="2012-01-01" gender="M" lastname="Schäfer" firstname="Conrad" license="445622">
              <RESULTS>
                <RESULT resultid="1002" eventid="6" swimtime="00:00:47.31" lane="2" heatid="6003" />
                <RESULT resultid="1001" eventid="11" swimtime="00:01:46.64" lane="2" heatid="11003" />
                <RESULT resultid="1000" eventid="13" swimtime="00:00:41.05" lane="8" heatid="13003" />
                <RESULT resultid="999" eventid="22" swimtime="00:00:54.50" lane="7" heatid="22009" />
                <RESULT resultid="998" eventid="24" swimtime="00:03:17.60" lane="3" heatid="24002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:37.50" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="997" eventid="32" swimtime="00:00:59.63" lane="3" heatid="32003" />
                <RESULT resultid="996" eventid="34" swimtime="00:01:31.52" lane="1" heatid="34002" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="189" birthdate="2015-01-01" gender="F" lastname="Beck" firstname="Charlotte" license="463336">
              <RESULTS>
                <RESULT resultid="1006" eventid="19" swimtime="00:01:01.39" lane="4" heatid="19005" />
                <RESULT resultid="1005" eventid="25" swimtime="00:01:00.85" lane="3" heatid="25003" />
                <RESULT resultid="1004" eventid="27" swimtime="00:01:11.40" lane="6" heatid="27004" />
                <RESULT resultid="1003" eventid="29" swimtime="00:01:01.11" lane="2" heatid="29003" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="190" birthdate="2014-01-01" gender="M" lastname="Al-Jumaili" firstname="Anas" license="446743">
              <RESULTS>
                <RESULT resultid="1010" eventid="20" swimtime="00:01:03.14" lane="7" heatid="20005" />
                <RESULT resultid="1009" eventid="26" swimtime="00:00:58.10" lane="1" heatid="26006" />
                <RESULT resultid="1008" eventid="28" swimtime="00:01:15.64" lane="3" heatid="28002" />
                <RESULT resultid="1007" eventid="30" swimtime="00:00:56.38" lane="2" heatid="30003" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="191" birthdate="2014-01-01" gender="M" lastname="Sommer" firstname="Alfred" license="446746">
              <RESULTS>
                <RESULT resultid="1015" eventid="18" status="WDR" swimtime="00:00:00.00" lane="4" heatid="18004" />
                <RESULT resultid="1014" eventid="22" status="WDR" swimtime="00:00:00.00" lane="4" heatid="22005" />
                <RESULT resultid="1013" eventid="26" status="WDR" swimtime="00:00:00.00" lane="8" heatid="26010" />
                <RESULT resultid="1012" eventid="30" status="WDR" swimtime="00:00:00.00" lane="3" heatid="30005" />
                <RESULT resultid="1011" eventid="34" status="WDR" swimtime="00:00:00.00" lane="5" heatid="34002" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="192" birthdate="2014-01-01" gender="M" lastname="Hache" firstname="Alexander" license="463410">
              <RESULTS>
                <RESULT resultid="1020" eventid="20" swimtime="00:00:53.21" lane="1" heatid="20011" />
                <RESULT resultid="1019" eventid="26" swimtime="00:00:44.86" lane="3" heatid="26015" />
                <RESULT resultid="1018" eventid="28" swimtime="00:00:58.71" lane="3" heatid="28007" />
                <RESULT resultid="1017" eventid="30" swimtime="00:00:40.63" lane="6" heatid="30008" />
                <RESULT resultid="1016" eventid="34" swimtime="00:01:34.01" lane="7" heatid="34004" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="ST Erzgebirge" nation="GER" region="12" code="5134">
          <ATHLETES>
            <ATHLETE athleteid="780" birthdate="2008-01-01" gender="M" lastname="Kulai" firstname="Vasyl" license="429668">
              <RESULTS>
                <RESULT resultid="3716" eventid="2" swimtime="00:03:08.04" lane="3" heatid="2001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:29.87" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="3715" eventid="15" swimtime="00:03:11.02" lane="6" heatid="15006">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:30.40" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="3714" eventid="20" swimtime="00:00:39.04" lane="7" heatid="20020" />
                <RESULT resultid="3713" eventid="34" swimtime="00:01:16.03" lane="3" heatid="34011" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="781" birthdate="2014-01-01" gender="F" lastname="Viertel" firstname="Victoria-Luise" license="461991">
              <RESULTS>
                <RESULT resultid="3719" eventid="19" swimtime="00:00:59.85" lane="2" heatid="19007" />
                <RESULT resultid="3718" eventid="25" swimtime="00:01:03.68" lane="6" heatid="25009" />
                <RESULT resultid="3717" eventid="27" swimtime="00:01:07.89" lane="3" heatid="27004" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="782" birthdate="2008-01-01" gender="F" lastname="Richter" firstname="Tine" license="429666">
              <RESULTS>
                <RESULT resultid="3724" eventid="1" swimtime="00:03:25.08" lane="3" heatid="1001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:32.10" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="3723" eventid="5" swimtime="00:00:38.61" lane="6" heatid="5008" />
                <RESULT resultid="3722" eventid="12" swimtime="00:00:32.31" lane="5" heatid="12015" />
                <RESULT resultid="3721" eventid="23" swimtime="00:02:55.05" lane="2" heatid="23001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:22.29" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="3720" eventid="35" swimtime="00:01:39.47" lane="2" heatid="35002" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="783" birthdate="2007-01-01" gender="F" lastname="Steiner" firstname="Tiffany" license="355425">
              <RESULTS>
                <RESULT resultid="3726" eventid="25" swimtime="00:00:37.08" lane="5" heatid="25032" />
                <RESULT resultid="3725" eventid="33" swimtime="00:01:13.48" lane="7" heatid="33016" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="784" birthdate="2013-01-01" gender="F" lastname="Oestreich" firstname="Sophia" license="458275">
              <RESULTS>
                <RESULT resultid="3731" eventid="10" swimtime="00:01:55.19" lane="3" heatid="10002" />
                <RESULT resultid="3730" eventid="12" swimtime="00:00:42.51" lane="5" heatid="12002" />
                <RESULT resultid="3729" eventid="21" swimtime="00:00:58.49" lane="6" heatid="21003" />
                <RESULT resultid="3728" eventid="25" swimtime="00:00:51.11" lane="8" heatid="25015" />
                <RESULT resultid="3727" eventid="33" swimtime="00:01:40.71" lane="1" heatid="33003" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="785" birthdate="2010-01-01" gender="M" lastname="Gläser" firstname="Simon" license="461951">
              <RESULTS>
                <RESULT resultid="3734" eventid="20" swimtime="00:00:46.35" lane="3" heatid="20015" />
                <RESULT resultid="3733" eventid="24" swimtime="00:03:11.37" lane="5" heatid="24001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:29.74" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="3732" eventid="34" swimtime="00:01:25.33" lane="3" heatid="34004" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="786" birthdate="2013-01-01" gender="M" lastname="Meyer" firstname="Sammy" license="458126">
              <RESULTS>
                <RESULT resultid="3738" eventid="18" swimtime="00:01:11.63" lane="3" heatid="18001" />
                <RESULT resultid="3737" eventid="22" swimtime="00:01:00.40" lane="1" heatid="22006" />
                <RESULT resultid="3736" eventid="26" swimtime="00:00:53.20" lane="2" heatid="26009" />
                <RESULT resultid="3735" eventid="34" swimtime="00:01:38.26" lane="4" heatid="34002" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="787" birthdate="2011-01-01" gender="F" lastname="Neubert" firstname="Sally" license="429664">
              <RESULTS>
                <RESULT resultid="3743" eventid="5" swimtime="00:00:54.60" lane="2" heatid="5003" />
                <RESULT resultid="3742" eventid="10" swimtime="00:01:49.91" lane="3" heatid="10003" />
                <RESULT resultid="3741" eventid="12" swimtime="00:00:43.22" lane="8" heatid="12003" />
                <RESULT resultid="3740" eventid="25" swimtime="00:00:51.37" lane="7" heatid="25016" />
                <RESULT resultid="3739" eventid="33" swimtime="00:01:35.03" lane="3" heatid="33004" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="788" birthdate="2007-01-01" gender="F" lastname="Hermann" firstname="Rebekka" license="402476">
              <RESULTS>
                <RESULT resultid="3745" eventid="23" swimtime="00:03:12.43" lane="7" heatid="23001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:26.40" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="3744" eventid="33" swimtime="00:01:19.24" lane="1" heatid="33009" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="789" birthdate="2012-01-01" gender="M" lastname="Bochmann" firstname="Noa" license="461952">
              <RESULTS>
                <RESULT resultid="3751" eventid="4" swimtime="00:01:57.65" lane="2" heatid="4002" />
                <RESULT resultid="3750" eventid="13" swimtime="00:00:46.73" lane="1" heatid="13002" />
                <RESULT resultid="3749" eventid="20" swimtime="00:00:54.65" lane="7" heatid="20007" />
                <RESULT resultid="3748" eventid="22" swimtime="00:01:07.39" lane="6" heatid="22002" />
                <RESULT resultid="3747" eventid="28" swimtime="00:01:07.11" lane="5" heatid="28002" />
                <RESULT resultid="3746" eventid="34" swimtime="00:01:45.76" lane="6" heatid="34001" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="790" birthdate="2010-01-01" gender="F" lastname="Lorenz" firstname="Milena" license="417871">
              <RESULTS>
                <RESULT resultid="3753" eventid="25" swimtime="00:00:52.80" lane="2" heatid="25016" />
                <RESULT resultid="3752" eventid="33" swimtime="00:01:39.78" lane="5" heatid="33005" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="791" birthdate="2012-01-01" gender="F" lastname="Langer" firstname="Mia" license="461959">
              <RESULTS>
                <RESULT resultid="3757" eventid="21" status="DNS" swimtime="00:00:00.00" lane="6" heatid="21007" />
                <RESULT resultid="3756" eventid="27" status="DNS" swimtime="00:00:00.00" lane="7" heatid="27002" />
                <RESULT resultid="3755" eventid="31" status="DNS" swimtime="00:00:00.00" lane="6" heatid="31002" />
                <RESULT resultid="3754" eventid="33" status="DNS" swimtime="00:00:00.00" lane="6" heatid="33003" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="792" birthdate="2011-01-01" gender="F" lastname="Schreiter" firstname="Melissa" license="447078">
              <RESULTS>
                <RESULT resultid="3764" eventid="3" status="DNS" swimtime="00:00:00.00" lane="5" heatid="3009" />
                <RESULT resultid="3763" eventid="5" status="DNS" swimtime="00:00:00.00" lane="6" heatid="5007" />
                <RESULT resultid="3762" eventid="10" swimtime="00:01:33.10" lane="7" heatid="10005" />
                <RESULT resultid="3761" eventid="14" swimtime="00:03:23.79" lane="1" heatid="14006">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:36.76" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="3760" eventid="19" swimtime="00:00:46.09" lane="8" heatid="19023" />
                <RESULT resultid="3759" eventid="23" swimtime="00:02:54.03" lane="7" heatid="23004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:23.76" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="3758" eventid="33" status="DNS" swimtime="00:00:00.00" lane="8" heatid="33009" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="793" birthdate="2013-01-01" gender="M" lastname="Nordheim" firstname="Matteo" license="461956">
              <RESULTS>
                <RESULT resultid="3767" eventid="18" status="DNS" swimtime="00:00:00.00" lane="4" heatid="18001" />
                <RESULT resultid="3766" eventid="22" status="DNS" swimtime="00:00:00.00" lane="1" heatid="22001" />
                <RESULT resultid="3765" eventid="32" status="DNS" swimtime="00:00:00.00" lane="5" heatid="32001" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="794" birthdate="2009-01-01" gender="M" lastname="Tutzschky" firstname="Lukas" license="461949">
              <RESULTS>
                <RESULT resultid="3771" eventid="6" swimtime="00:00:40.30" lane="6" heatid="6006" />
                <RESULT resultid="3770" eventid="13" swimtime="00:00:33.76" lane="4" heatid="13008" />
                <RESULT resultid="3769" eventid="24" swimtime="00:02:55.27" lane="4" heatid="24003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:24.26" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="3768" eventid="34" swimtime="00:01:18.47" lane="7" heatid="34007" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="795" birthdate="2010-01-01" gender="F" lastname="Göhler" firstname="Lucy" license="402479">
              <RESULTS>
                <RESULT resultid="3773" eventid="23" swimtime="00:02:51.33" lane="7" heatid="23006">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:22.84" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="3772" eventid="33" swimtime="00:01:18.26" lane="6" heatid="33010" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="796" birthdate="2008-01-01" gender="M" lastname="Heidenreich" firstname="Luca" license="415867">
              <RESULTS>
                <RESULT resultid="3778" eventid="4" swimtime="00:01:22.11" lane="6" heatid="4011" />
                <RESULT resultid="3777" eventid="6" swimtime="00:00:34.91" lane="7" heatid="6008" />
                <RESULT resultid="3776" eventid="15" swimtime="00:02:58.49" lane="3" heatid="15007">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:27.17" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="3775" eventid="20" swimtime="00:00:34.95" lane="2" heatid="20022" />
                <RESULT resultid="3774" eventid="26" swimtime="00:00:36.15" lane="1" heatid="26023" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="797" birthdate="2011-01-01" gender="F" lastname="Rößler" firstname="Lina" license="476556">
              <RESULTS>
                <RESULT resultid="3782" eventid="5" status="DSQ" swimtime="00:00:58.52" lane="2" heatid="5001" comment="Letzter Armzug nicht über Wasser nach vorn gebracht." />
                <RESULT resultid="3781" eventid="10" swimtime="00:02:06.74" lane="3" heatid="10001" />
                <RESULT resultid="3780" eventid="19" swimtime="00:00:58.88" lane="7" heatid="19001" />
                <RESULT resultid="3779" eventid="25" swimtime="00:00:53.97" lane="3" heatid="25001" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="798" birthdate="2007-01-01" gender="M" lastname="Richter" firstname="Kimi" license="384061">
              <RESULTS>
                <RESULT resultid="3786" eventid="11" status="DNS" swimtime="00:00:00.00" lane="6" heatid="11012" />
                <RESULT resultid="3785" eventid="13" status="DNS" swimtime="00:00:00.00" lane="5" heatid="13017" />
                <RESULT resultid="3784" eventid="26" swimtime="00:00:30.76" lane="3" heatid="26024" />
                <RESULT resultid="3783" eventid="38" swimtime="00:02:34.45" lane="2" heatid="38005">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:14.94" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="799" birthdate="2012-01-01" gender="M" lastname="Gottschalk" firstname="Karl" license="461957">
              <RESULTS>
                <RESULT resultid="3791" eventid="4" status="DSQ" swimtime="00:01:56.24" lane="5" heatid="4002" comment="Start vor dem Startsignal." />
                <RESULT resultid="3790" eventid="13" swimtime="00:00:45.45" lane="3" heatid="13001" />
                <RESULT resultid="3789" eventid="20" swimtime="00:00:53.21" lane="1" heatid="20016" />
                <RESULT resultid="3788" eventid="22" status="DSQ" swimtime="00:01:17.70" lane="2" heatid="22001" comment="Das Brett wurde beim Zielanschlag nicht am vorderen Rand umfasst." />
                <RESULT resultid="3787" eventid="28" swimtime="00:01:05.29" lane="2" heatid="28004" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="800" birthdate="2014-01-01" gender="M" lastname="Gläser" firstname="Julian" license="458122">
              <RESULTS>
                <RESULT resultid="3795" eventid="18" status="DNS" swimtime="00:00:00.00" lane="4" heatid="18006" />
                <RESULT resultid="3794" eventid="22" status="DNS" swimtime="00:00:00.00" lane="4" heatid="22008" />
                <RESULT resultid="3793" eventid="30" status="DNS" swimtime="00:00:00.00" lane="8" heatid="30005" />
                <RESULT resultid="3792" eventid="34" status="DNS" swimtime="00:00:00.00" lane="2" heatid="34001" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="801" birthdate="2007-01-01" gender="M" lastname="Neubert" firstname="Johannes" license="393375">
              <RESULTS>
                <RESULT resultid="3799" eventid="4" swimtime="00:01:27.08" lane="3" heatid="4009" />
                <RESULT resultid="3798" eventid="13" swimtime="00:00:30.34" lane="2" heatid="13015" />
                <RESULT resultid="3797" eventid="20" swimtime="00:00:38.36" lane="2" heatid="20020" />
                <RESULT resultid="3796" eventid="34" swimtime="00:01:09.53" lane="5" heatid="34012" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="802" birthdate="2013-01-01" gender="M" lastname="Lehmann" firstname="Jay" license="461955">
              <RESULTS>
                <RESULT resultid="3804" eventid="6" swimtime="00:00:58.59" lane="1" heatid="6001" />
                <RESULT resultid="3803" eventid="13" swimtime="00:00:48.48" lane="4" heatid="13001" />
                <RESULT resultid="3802" eventid="22" status="DSQ" swimtime="00:01:14.07" lane="7" heatid="22001" comment="Das Brett wurde beim Zielanschlag nicht umfasst." />
                <RESULT resultid="3801" eventid="32" swimtime="00:01:17.06" lane="3" heatid="32001" />
                <RESULT resultid="3800" eventid="34" swimtime="00:01:43.14" lane="5" heatid="34001" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="803" birthdate="2013-01-01" gender="M" lastname="Rebentrost" firstname="Helios" license="461954">
              <RESULTS>
                <RESULT resultid="3807" eventid="6" swimtime="00:00:53.00" lane="5" heatid="6001" />
                <RESULT resultid="3806" eventid="11" swimtime="00:01:54.66" lane="1" heatid="11002" />
                <RESULT resultid="3805" eventid="13" swimtime="00:00:50.24" lane="8" heatid="13002" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="804" birthdate="2007-01-01" gender="F" lastname="Schönherr" firstname="Hannah" license="382221">
              <RESULTS>
                <RESULT resultid="3809" eventid="25" swimtime="00:00:44.23" lane="8" heatid="25028" />
                <RESULT resultid="3808" eventid="35" swimtime="00:01:52.26" lane="6" heatid="35002" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="805" birthdate="2012-01-01" gender="F" lastname="Müller" firstname="Frieda" license="461992">
              <RESULTS>
                <RESULT resultid="3812" eventid="19" swimtime="00:00:51.88" lane="7" heatid="19015" />
                <RESULT resultid="3811" eventid="25" swimtime="00:00:46.52" lane="4" heatid="25016" />
                <RESULT resultid="3810" eventid="33" swimtime="00:01:28.61" lane="8" heatid="33006" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="806" birthdate="2011-01-01" gender="M" lastname="Fauska" firstname="Franz" license="458123">
              <RESULTS>
                <RESULT resultid="3815" eventid="4" swimtime="00:01:51.14" lane="3" heatid="4003" />
                <RESULT resultid="3814" eventid="13" swimtime="00:00:42.52" lane="6" heatid="13002" />
                <RESULT resultid="3813" eventid="15" swimtime="00:03:59.28" lane="2" heatid="15002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:58.71" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="807" birthdate="2009-01-01" gender="M" lastname="Findeisen" firstname="Erik" license="415866">
              <RESULTS>
                <RESULT resultid="3819" eventid="6" status="DNS" swimtime="00:00:00.00" lane="4" heatid="6009" />
                <RESULT resultid="3818" eventid="13" status="DNS" swimtime="00:00:00.00" lane="7" heatid="13016" />
                <RESULT resultid="3817" eventid="20" swimtime="00:00:38.20" lane="7" heatid="20021" />
                <RESULT resultid="3816" eventid="36" swimtime="00:01:20.41" lane="4" heatid="36002" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="808" birthdate="2009-01-01" gender="F" lastname="Wittig" firstname="Emma" license="415865">
              <RESULTS>
                <RESULT resultid="3823" eventid="3" swimtime="00:01:24.50" lane="6" heatid="3011" />
                <RESULT resultid="3822" eventid="14" swimtime="00:03:14.10" lane="7" heatid="14007">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:32.32" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="3821" eventid="19" swimtime="00:00:37.74" lane="5" heatid="19026" />
                <RESULT resultid="3820" eventid="35" swimtime="00:01:24.29" lane="6" heatid="35003" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="809" birthdate="2013-01-01" gender="F" lastname="Klaus" firstname="Emma" license="461960">
              <RESULTS>
                <RESULT resultid="3828" eventid="3" swimtime="00:01:56.91" lane="5" heatid="3002" />
                <RESULT resultid="3827" eventid="14" swimtime="00:04:12.42" lane="3" heatid="14001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:02:01.52" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="3826" eventid="19" swimtime="00:00:53.76" lane="7" heatid="19014" />
                <RESULT resultid="3825" eventid="27" swimtime="00:01:04.21" lane="7" heatid="27009" />
                <RESULT resultid="3824" eventid="31" swimtime="00:01:20.98" lane="8" heatid="31002" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="810" birthdate="2015-01-01" gender="F" lastname="Morgenstern" firstname="Elena" license="471532">
              <RESULTS>
                <RESULT resultid="3832" eventid="19" swimtime="00:00:55.99" lane="1" heatid="19007" />
                <RESULT resultid="3831" eventid="25" swimtime="00:00:56.92" lane="4" heatid="25006" />
                <RESULT resultid="3830" eventid="27" swimtime="00:01:05.89" lane="4" heatid="27001" />
                <RESULT resultid="3829" eventid="29" swimtime="00:01:00.00" lane="5" heatid="29002" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="811" birthdate="2009-01-01" gender="M" lastname="Neubert" firstname="Domenic" license="429667">
              <RESULTS>
                <RESULT resultid="3836" eventid="2" swimtime="00:03:11.30" lane="5" heatid="2001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:32.12" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="3835" eventid="11" swimtime="00:01:31.11" lane="6" heatid="11008" />
                <RESULT resultid="3834" eventid="26" swimtime="00:00:39.73" lane="2" heatid="26021" />
                <RESULT resultid="3833" eventid="36" status="DSQ" swimtime="00:01:35.64" lane="6" heatid="36002" comment="Der Sportler führte auf der Schwimmstrecke mehrere Wechselbeinschläge aus." />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="812" birthdate="2013-01-01" gender="M" lastname="Konrad" firstname="Christian" license="461953">
              <RESULTS>
                <RESULT resultid="3840" eventid="20" swimtime="00:00:52.00" lane="1" heatid="20010" />
                <RESULT resultid="3839" eventid="22" swimtime="00:00:59.23" lane="1" heatid="22005" />
                <RESULT resultid="3838" eventid="28" swimtime="00:01:08.04" lane="5" heatid="28001" />
                <RESULT resultid="3837" eventid="32" swimtime="00:01:07.16" lane="4" heatid="32003" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="813" birthdate="2015-01-01" gender="M" lastname="Unger" firstname="Bruno" license="471531">
              <RESULTS>
                <RESULT resultid="3844" eventid="20" swimtime="00:00:55.33" lane="7" heatid="20009" />
                <RESULT resultid="3843" eventid="22" swimtime="00:01:11.97" lane="3" heatid="22005" />
                <RESULT resultid="3842" eventid="28" swimtime="00:01:01.36" lane="8" heatid="28005" />
                <RESULT resultid="3841" eventid="30" swimtime="00:00:54.17" lane="8" heatid="30003" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="814" birthdate="2011-01-01" gender="F" lastname="Müller" firstname="Annica" license="429663">
              <RESULTS>
                <RESULT resultid="3846" eventid="23" swimtime="00:02:48.48" lane="6" heatid="23006">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:21.61" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="3845" eventid="33" swimtime="00:01:13.00" lane="3" heatid="33012" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="815" birthdate="2010-01-01" gender="M" lastname="Neubert" firstname="Alois" license="461950">
              <RESULTS>
                <RESULT resultid="3850" eventid="4" swimtime="00:02:09.70" lane="4" heatid="4001" />
                <RESULT resultid="3849" eventid="13" swimtime="00:00:44.56" lane="5" heatid="13002" />
                <RESULT resultid="3848" eventid="20" swimtime="00:00:58.59" lane="6" heatid="20006" />
                <RESULT resultid="3847" eventid="26" swimtime="00:00:52.91" lane="2" heatid="26008" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1379" birthdate="2011-01-01" gender="F" lastname="Hiemann" firstname="Elisa" license="447078">
              <RESULTS>
                <RESULT resultid="6359" eventid="3" swimtime="00:01:37.11" lane="6" heatid="3001" />
                <RESULT resultid="6362" eventid="5" swimtime="00:00:44.17" lane="7" heatid="5001" />
                <RESULT resultid="6361" eventid="14" swimtime="00:03:39.71" lane="2" heatid="14001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:51.31" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="6360" eventid="19" swimtime="00:00:43.43" lane="8" heatid="19001" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY number="1" gender="X" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="3851" eventid="7" swimtime="00:03:02.52" lane="4" heatid="7001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:28.19" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="792" number="1" />
                    <RELAYPOSITION athleteid="1379" number="2" />
                    <RELAYPOSITION athleteid="803" number="3" />
                    <RELAYPOSITION athleteid="815" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" gender="X" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="6366" eventid="16" status="DNS" swimtime="00:00:00.00" lane="3" heatid="16001" />
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB name="Startgemeinschaft Dresden" nation="GER" region="20" code="0">
          <ATHLETES>
            <ATHLETE athleteid="843" birthdate="2009-01-01" gender="F" lastname="Zimmermanns" firstname="Ariane" license="0">
              <RESULTS>
                <RESULT resultid="3970" eventid="41" status="DSQ" swimtime="00:00:23.44" lane="5" heatid="41001" comment="Gesicht aus dem Wasser." />
                <RESULT resultid="3971" eventid="45" swimtime="00:01:14.45" lane="7" heatid="45003" />
                <RESULT resultid="3972" eventid="49" status="DNS" swimtime="00:00:00.00" lane="3" heatid="49002" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="844" birthdate="2009-01-01" gender="M" lastname="Hübner" firstname="Christoph" license="0">
              <RESULTS>
                <RESULT resultid="3973" eventid="42" status="DSQ" swimtime="00:00:18.91" lane="5" heatid="42002" comment="Gesicht aus dem Wasser." />
                <RESULT resultid="3974" eventid="46" swimtime="00:01:11.86" lane="6" heatid="46002" />
                <RESULT resultid="3975" eventid="50" swimtime="00:00:29.80" lane="8" heatid="50003" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="845" birthdate="2012-01-01" gender="F" lastname="Körner" firstname="Ella Henriette" license="0">
              <RESULTS>
                <RESULT resultid="3976" eventid="41" swimtime="00:00:16.22" lane="2" heatid="41002" />
                <RESULT resultid="3977" eventid="45" swimtime="00:01:12.36" lane="2" heatid="45004" />
                <RESULT resultid="3978" eventid="49" swimtime="00:00:32.09" lane="7" heatid="49003" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="846" birthdate="2012-01-01" gender="F" lastname="Bernhardt" firstname="Fjora" license="0">
              <RESULTS>
                <RESULT resultid="3979" eventid="41" swimtime="00:00:19.50" lane="4" heatid="41001" />
                <RESULT resultid="3980" eventid="45" swimtime="00:01:15.62" lane="1" heatid="45003" />
                <RESULT resultid="3981" eventid="49" swimtime="00:00:33.44" lane="7" heatid="49002" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="847" birthdate="2013-01-01" gender="M" lastname="Schewitzer" firstname="Gustav" license="0">
              <RESULTS>
                <RESULT resultid="3982" eventid="42" swimtime="00:00:17.03" lane="1" heatid="42003" />
                <RESULT resultid="3983" eventid="46" swimtime="00:01:13.03" lane="1" heatid="46003" />
                <RESULT resultid="3984" eventid="50" status="DSQ" swimtime="00:00:31.32" lane="6" heatid="50003" comment="Falscher Start." />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="848" birthdate="2010-01-01" gender="F" lastname="Mucha" firstname="Helene" license="0">
              <RESULTS>
                <RESULT resultid="3985" eventid="41" swimtime="00:00:17.77" lane="1" heatid="41002" />
                <RESULT resultid="3986" eventid="45" swimtime="00:01:10.63" lane="3" heatid="45003" />
                <RESULT resultid="3987" eventid="49" swimtime="00:00:31.85" lane="4" heatid="49002" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="849" birthdate="2006-01-01" gender="F" lastname="Neumann" firstname="Josephine" license="0">
              <RESULTS>
                <RESULT resultid="3988" eventid="41" swimtime="00:00:13.26" lane="1" heatid="41005" />
                <RESULT resultid="3989" eventid="45" swimtime="00:01:01.32" lane="8" heatid="45006" />
                <RESULT resultid="3990" eventid="49" status="DNS" swimtime="00:00:00.00" lane="3" heatid="49004" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="850" birthdate="2006-01-01" gender="F" lastname="Schürer" firstname="Katka" license="0">
              <RESULTS>
                <RESULT resultid="3991" eventid="41" status="DSQ" swimtime="00:00:17.34" lane="5" heatid="41003" comment="zu zeitig aufgetaucht, vor Zielanschlag." />
                <RESULT resultid="3992" eventid="45" swimtime="00:01:10.48" lane="8" heatid="45005" />
                <RESULT resultid="3993" eventid="49" swimtime="00:00:30.61" lane="5" heatid="49003" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="851" birthdate="2010-01-01" gender="F" lastname="Kirchner" firstname="Klara" license="0">
              <RESULTS>
                <RESULT resultid="3994" eventid="41" status="DNS" swimtime="00:00:00.00" lane="8" heatid="41002" />
                <RESULT resultid="3995" eventid="45" status="DNS" swimtime="00:00:00.00" lane="5" heatid="45003" />
                <RESULT resultid="3996" eventid="49" status="DNS" swimtime="00:00:00.00" lane="2" heatid="49003" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="852" birthdate="2007-01-01" gender="F" lastname="Marquardt" firstname="Lotte" license="0">
              <RESULTS>
                <RESULT resultid="3997" eventid="39" swimtime="00:02:12.01" lane="7" heatid="39003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:02.96" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="3998" eventid="41" swimtime="00:00:13.05" lane="2" heatid="41005" />
                <RESULT resultid="3999" eventid="45" swimtime="00:01:01.06" lane="7" heatid="45006" />
                <RESULT resultid="4000" eventid="49" swimtime="00:00:27.97" lane="8" heatid="49005" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="853" birthdate="2007-01-01" gender="F" lastname="Bretschneider" firstname="Luisa" license="0">
              <RESULTS>
                <RESULT resultid="4001" eventid="39" swimtime="00:02:35.17" lane="8" heatid="39002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:14.04" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="4002" eventid="41" swimtime="00:00:14.67" lane="4" heatid="41003" />
                <RESULT resultid="4003" eventid="45" swimtime="00:01:08.80" lane="1" heatid="45004" />
                <RESULT resultid="4004" eventid="49" swimtime="00:00:29.86" lane="4" heatid="49003" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="854" birthdate="2011-01-01" gender="M" lastname="Buchmann" firstname="Marco" license="0">
              <RESULTS>
                <RESULT resultid="4005" eventid="42" swimtime="00:00:17.52" lane="3" heatid="42002" />
                <RESULT resultid="4006" eventid="46" swimtime="00:01:10.93" lane="3" heatid="46002" />
                <RESULT resultid="4007" eventid="50" swimtime="00:00:31.17" lane="7" heatid="50003" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="855" birthdate="2011-01-01" gender="F" lastname="Gey" firstname="Mathilde" license="0">
              <RESULTS>
                <RESULT resultid="4008" eventid="41" swimtime="00:00:19.09" lane="7" heatid="41003" />
                <RESULT resultid="4009" eventid="45" swimtime="00:01:12.23" lane="5" heatid="45004" />
                <RESULT resultid="4010" eventid="49" swimtime="00:00:32.34" lane="3" heatid="49003" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="856" birthdate="2011-01-01" gender="F" lastname="Oehme" firstname="Mia" license="0">
              <RESULTS>
                <RESULT resultid="4011" eventid="41" swimtime="00:00:18.02" lane="7" heatid="41002" />
                <RESULT resultid="4012" eventid="45" swimtime="00:01:11.86" lane="8" heatid="45004" />
                <RESULT resultid="4013" eventid="49" status="DSQ" swimtime="00:00:00.00" lane="8" heatid="49003" comment="Aufgegeben." />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="857" birthdate="2011-01-01" gender="F" lastname="Müller" firstname="Reni" license="0">
              <RESULTS>
                <RESULT resultid="4014" eventid="41" swimtime="00:00:17.36" lane="1" heatid="41003" />
                <RESULT resultid="4015" eventid="45" swimtime="00:01:11.19" lane="4" heatid="45004" />
                <RESULT resultid="4016" eventid="49" swimtime="00:00:31.91" lane="6" heatid="49003" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="858" birthdate="2007-01-01" gender="F" lastname="Razumovska" firstname="Sophiya" license="0">
              <RESULTS>
                <RESULT resultid="4017" eventid="41" status="DSQ" swimtime="00:00:12.88" lane="5" heatid="41004" comment="Becken über die Anschlagmatte verlassen." />
                <RESULT resultid="4018" eventid="45" swimtime="00:01:03.56" lane="6" heatid="45005" />
                <RESULT resultid="4019" eventid="49" swimtime="00:00:26.62" lane="4" heatid="49004" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="STV Limbach-Oberfrohna e.V." nation="GER" region="12" code="5406">
          <ATHLETES>
            <ATHLETE athleteid="1052" birthdate="2012-01-01" gender="F" lastname="Lienert" firstname="Alexa" license="408032">
              <RESULTS>
                <RESULT resultid="4917" eventid="5" swimtime="00:00:43.39" lane="1" heatid="5005" />
                <RESULT resultid="4918" eventid="10" swimtime="00:01:36.28" lane="4" heatid="10003" />
                <RESULT resultid="4919" eventid="12" swimtime="00:00:37.86" lane="4" heatid="12007" />
                <RESULT resultid="4920" eventid="19" swimtime="00:00:52.33" lane="3" heatid="19013" />
                <RESULT resultid="4921" eventid="25" swimtime="00:00:44.85" lane="3" heatid="25022" />
                <RESULT resultid="4922" eventid="35" swimtime="00:01:45.72" lane="7" heatid="35002" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1053" birthdate="2015-01-01" gender="M" lastname="Ronneburger" firstname="Collin" license="460545">
              <RESULTS>
                <RESULT resultid="4923" eventid="20" status="DSQ" swimtime="00:01:05.01" lane="1" heatid="20006" comment="Vor dem Ziel wurden die Hände weiter als bis zur Hüftlinie nach hinten gebracht." />
                <RESULT resultid="4924" eventid="28" swimtime="00:01:05.12" lane="2" heatid="28005" />
                <RESULT resultid="4925" eventid="30" swimtime="00:00:49.51" lane="5" heatid="30006" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1054" birthdate="2011-01-01" gender="F" lastname="Türk" firstname="Emilia" license="408039">
              <RESULTS>
                <RESULT resultid="4926" eventid="1" swimtime="00:03:10.67" lane="4" heatid="1003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:29.70" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="4927" eventid="5" swimtime="00:00:42.73" lane="8" heatid="5006" />
                <RESULT resultid="4928" eventid="10" swimtime="00:01:29.51" lane="2" heatid="10008" />
                <RESULT resultid="4929" eventid="12" swimtime="00:00:34.74" lane="3" heatid="12011" />
                <RESULT resultid="4930" eventid="23" swimtime="00:02:47.70" lane="1" heatid="23008">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:21.10" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="4931" eventid="25" swimtime="00:00:42.62" lane="7" heatid="25028" />
                <RESULT resultid="4932" eventid="33" swimtime="00:01:16.31" lane="4" heatid="33010" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1055" birthdate="2010-01-01" gender="F" lastname="Reschke" firstname="Fanny Florentine" license="421222">
              <RESULTS>
                <RESULT resultid="4933" eventid="23" swimtime="00:02:46.41" lane="8" heatid="23010">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:18.85" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="4934" eventid="25" swimtime="00:00:40.01" lane="3" heatid="25030" />
                <RESULT resultid="4935" eventid="33" swimtime="00:01:14.85" lane="7" heatid="33014" />
                <RESULT resultid="4936" eventid="37" swimtime="00:03:07.39" lane="8" heatid="37007">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:32.82" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1056" birthdate="2015-01-01" gender="F" lastname="Ettelt" firstname="Hanna" license="471930">
              <RESULTS>
                <RESULT resultid="4937" eventid="19" swimtime="00:01:03.78" lane="2" heatid="19004" />
                <RESULT resultid="4938" eventid="25" swimtime="00:01:10.65" lane="1" heatid="25002" />
                <RESULT resultid="4939" eventid="27" swimtime="00:01:24.45" lane="2" heatid="27002" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1057" birthdate="2009-01-01" gender="F" lastname="Lienert" firstname="Mareike" license="387936">
              <RESULTS>
                <RESULT resultid="4940" eventid="5" swimtime="00:00:33.14" lane="8" heatid="5013" />
                <RESULT resultid="4941" eventid="10" swimtime="00:01:20.25" lane="7" heatid="10014" />
                <RESULT resultid="4942" eventid="12" swimtime="00:00:30.50" lane="5" heatid="12017" />
                <RESULT resultid="4943" eventid="19" swimtime="00:00:43.03" lane="2" heatid="19025" />
                <RESULT resultid="4944" eventid="25" swimtime="00:00:37.37" lane="2" heatid="25033" />
                <RESULT resultid="4945" eventid="33" swimtime="00:01:11.87" lane="1" heatid="33017" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1058" birthdate="2012-01-01" gender="M" lastname="Hennig" firstname="Max" license="457928">
              <RESULTS>
                <RESULT resultid="4946" eventid="6" status="WDR" swimtime="00:00:00.00" lane="1" heatid="6003" />
                <RESULT resultid="4947" eventid="11" status="WDR" swimtime="00:00:00.00" lane="4" heatid="11003" />
                <RESULT resultid="4948" eventid="13" status="WDR" swimtime="00:00:00.00" lane="3" heatid="13005" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1059" birthdate="2008-01-01" gender="M" lastname="Rauchfuß" firstname="Max" license="393450">
              <RESULTS>
                <RESULT resultid="4949" eventid="4" swimtime="00:01:24.03" lane="2" heatid="4010" />
                <RESULT resultid="4950" eventid="6" swimtime="00:00:31.07" lane="7" heatid="6010" />
                <RESULT resultid="4951" eventid="13" swimtime="00:00:28.83" lane="3" heatid="13016" />
                <RESULT resultid="4952" eventid="15" swimtime="00:03:06.90" lane="3" heatid="15006">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:32.05" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="4953" eventid="20" swimtime="00:00:36.66" lane="1" heatid="20021" />
                <RESULT resultid="4954" eventid="34" swimtime="00:01:05.65" lane="8" heatid="34014" />
                <RESULT resultid="4955" eventid="36" swimtime="00:01:14.27" lane="2" heatid="36003" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1060" birthdate="2013-01-01" gender="F" lastname="Veit" firstname="Mia Sophie" license="451368">
              <RESULTS>
                <RESULT resultid="4956" eventid="3" swimtime="00:02:12.15" lane="7" heatid="3002" />
                <RESULT resultid="4957" eventid="5" swimtime="00:01:00.43" lane="6" heatid="5001" />
                <RESULT resultid="4958" eventid="10" swimtime="00:01:54.46" lane="2" heatid="10003" />
                <RESULT resultid="4959" eventid="12" swimtime="00:00:42.45" lane="3" heatid="12003" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="SV 1919 Grimma" nation="GER" region="12" code="5149">
          <ATHLETES>
            <ATHLETE athleteid="1068" birthdate="2013-01-01" gender="M" lastname="Munari" firstname="Alessandro" license="445022">
              <RESULTS>
                <RESULT resultid="4981" eventid="4" swimtime="00:01:59.30" lane="1" heatid="4003" />
                <RESULT resultid="4982" eventid="11" swimtime="00:01:31.98" lane="7" heatid="11007" />
                <RESULT resultid="4983" eventid="13" swimtime="00:00:38.27" lane="7" heatid="13005" />
                <RESULT resultid="4984" eventid="22" swimtime="00:00:51.05" lane="6" heatid="22010" />
                <RESULT resultid="4985" eventid="24" swimtime="00:03:02.18" lane="2" heatid="24005">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:27.39" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="4986" eventid="26" swimtime="00:00:43.15" lane="2" heatid="26016" />
                <RESULT resultid="4987" eventid="34" swimtime="00:01:23.48" lane="2" heatid="34007" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1069" birthdate="2010-01-01" gender="M" lastname="Duckstein" firstname="Alex" license="412300">
              <RESULTS>
                <RESULT resultid="4988" eventid="20" swimtime="00:00:47.10" lane="7" heatid="20014" />
                <RESULT resultid="4989" eventid="24" swimtime="00:02:57.34" lane="5" heatid="24004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:23.92" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="4990" eventid="26" swimtime="00:00:41.86" lane="4" heatid="26018" />
                <RESULT resultid="4991" eventid="34" swimtime="00:01:18.99" lane="6" heatid="34009" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1070" birthdate="2009-01-01" gender="F" lastname="Maneck" firstname="Amilia" license="398061">
              <RESULTS>
                <RESULT resultid="4992" eventid="1" swimtime="00:02:55.35" lane="2" heatid="1006">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:21.38" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="4993" eventid="5" swimtime="00:00:34.87" lane="5" heatid="5012" />
                <RESULT resultid="4994" eventid="10" swimtime="00:01:17.99" lane="6" heatid="10015" />
                <RESULT resultid="4995" eventid="12" swimtime="00:00:31.12" lane="2" heatid="12017" />
                <RESULT resultid="4996" eventid="25" swimtime="00:00:35.28" lane="6" heatid="25034" />
                <RESULT resultid="4997" eventid="33" swimtime="00:01:07.47" lane="7" heatid="33018" />
                <RESULT resultid="4998" eventid="35" swimtime="00:01:25.06" lane="5" heatid="35003" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1071" birthdate="2010-01-01" gender="F" lastname="Hartwig" firstname="Annika" license="471349">
              <RESULTS>
                <RESULT resultid="4999" eventid="3" swimtime="00:01:44.14" lane="8" heatid="3007" />
                <RESULT resultid="5000" eventid="5" swimtime="00:00:52.60" lane="1" heatid="5002" />
                <RESULT resultid="5001" eventid="12" swimtime="00:00:39.74" lane="7" heatid="12004" />
                <RESULT resultid="5002" eventid="19" swimtime="00:00:48.58" lane="1" heatid="19018" />
                <RESULT resultid="5003" eventid="25" swimtime="00:00:49.71" lane="3" heatid="25013" />
                <RESULT resultid="5004" eventid="33" swimtime="00:01:31.04" lane="2" heatid="33006" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1072" birthdate="2015-01-01" gender="F" lastname="Golze" firstname="Clara" license="463479">
              <RESULTS>
                <RESULT resultid="5005" eventid="17" swimtime="00:01:05.72" lane="1" heatid="17009" />
                <RESULT resultid="5006" eventid="19" swimtime="00:01:11.73" lane="4" heatid="19001" />
                <RESULT resultid="5007" eventid="25" swimtime="00:00:59.29" lane="6" heatid="25006" />
                <RESULT resultid="5008" eventid="27" swimtime="00:01:19.25" lane="4" heatid="27002" />
                <RESULT resultid="5009" eventid="29" swimtime="00:00:57.99" lane="5" heatid="29004" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1073" birthdate="2007-01-01" gender="F" lastname="Kösters" firstname="Constanze" license="393103">
              <RESULTS>
                <RESULT resultid="5010" eventid="5" swimtime="00:00:36.81" lane="1" heatid="5010" />
                <RESULT resultid="5011" eventid="8" swimtime="00:03:12.50" lane="5" heatid="8001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:27.99" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="5012" eventid="10" swimtime="00:01:19.67" lane="1" heatid="10015" />
                <RESULT resultid="5013" eventid="12" swimtime="00:00:34.90" lane="8" heatid="12012" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1074" birthdate="2015-01-01" gender="M" lastname="Schewelew" firstname="Egor" license="463483">
              <RESULTS>
                <RESULT resultid="5014" eventid="18" swimtime="00:01:12.66" lane="6" heatid="18004" />
                <RESULT resultid="5015" eventid="20" swimtime="00:01:02.07" lane="6" heatid="20003" />
                <RESULT resultid="5016" eventid="22" swimtime="00:01:18.79" lane="4" heatid="22001" />
                <RESULT resultid="5017" eventid="26" swimtime="00:00:50.88" lane="5" heatid="26006" />
                <RESULT resultid="5018" eventid="30" swimtime="00:00:47.15" lane="2" heatid="30006" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1075" birthdate="2014-01-01" gender="F" lastname="Brauße" firstname="Elena" license="451463">
              <RESULTS>
                <RESULT resultid="5019" eventid="19" swimtime="00:00:58.58" lane="4" heatid="19007" />
                <RESULT resultid="5020" eventid="25" swimtime="00:00:59.02" lane="7" heatid="25006" />
                <RESULT resultid="5021" eventid="27" status="DSQ" swimtime="00:01:06.65" lane="7" heatid="27007" comment="Wechselbeinschläge nach dem Start." />
                <RESULT resultid="5022" eventid="29" swimtime="00:00:51.05" lane="2" heatid="29004" />
                <RESULT resultid="5023" eventid="33" swimtime="00:02:01.08" lane="2" heatid="33002" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1076" birthdate="2014-01-01" gender="F" lastname="Streubel" firstname="Eliana Malea" license="451402">
              <RESULTS>
                <RESULT resultid="5024" eventid="19" swimtime="00:00:58.99" lane="5" heatid="19008" />
                <RESULT resultid="5025" eventid="21" swimtime="00:01:04.52" lane="8" heatid="21006" />
                <RESULT resultid="5026" eventid="27" swimtime="00:01:06.86" lane="7" heatid="27008" />
                <RESULT resultid="5027" eventid="29" swimtime="00:00:46.68" lane="1" heatid="29008" />
                <RESULT resultid="5028" eventid="33" swimtime="00:01:48.82" lane="3" heatid="33002" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1077" birthdate="2011-01-01" gender="F" lastname="Förster" firstname="Emily" license="436849">
              <RESULTS>
                <RESULT resultid="5029" eventid="19" swimtime="00:00:47.39" lane="3" heatid="19018" />
                <RESULT resultid="5030" eventid="23" swimtime="00:02:52.00" lane="3" heatid="23008">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:22.27" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="5031" eventid="25" swimtime="00:00:42.39" lane="6" heatid="25028" />
                <RESULT resultid="5032" eventid="33" swimtime="00:01:17.73" lane="5" heatid="33012" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1078" birthdate="2012-01-01" gender="F" lastname="Möbius" firstname="Emma" license="436843">
              <RESULTS>
                <RESULT resultid="5033" eventid="3" swimtime="00:01:48.26" lane="3" heatid="3004" />
                <RESULT resultid="5034" eventid="5" swimtime="00:00:49.96" lane="7" heatid="5003" />
                <RESULT resultid="5035" eventid="12" swimtime="00:00:38.57" lane="7" heatid="12006" />
                <RESULT resultid="5036" eventid="19" swimtime="00:00:50.13" lane="7" heatid="19018" />
                <RESULT resultid="5037" eventid="25" swimtime="00:00:44.21" lane="7" heatid="25021" />
                <RESULT resultid="5038" eventid="27" swimtime="00:00:56.52" lane="8" heatid="27012" />
                <RESULT resultid="5039" eventid="33" swimtime="00:01:30.44" lane="1" heatid="33007" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1079" birthdate="2015-01-01" gender="F" lastname="Päßler" firstname="Emma" license="463482">
              <RESULTS>
                <RESULT resultid="5040" eventid="17" swimtime="00:01:21.55" lane="8" heatid="17002" />
                <RESULT resultid="5041" eventid="21" swimtime="00:01:23.36" lane="8" heatid="21003" />
                <RESULT resultid="5042" eventid="25" swimtime="00:01:03.69" lane="2" heatid="25004" />
                <RESULT resultid="5043" eventid="29" swimtime="00:00:53.64" lane="6" heatid="29005" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1080" birthdate="2014-01-01" gender="F" lastname="Seemann" firstname="Emma" license="451406">
              <RESULTS>
                <RESULT resultid="5044" eventid="19" swimtime="00:00:55.97" lane="4" heatid="19011" />
                <RESULT resultid="5045" eventid="27" swimtime="00:01:08.37" lane="4" heatid="27006" />
                <RESULT resultid="5046" eventid="29" swimtime="00:00:44.77" lane="4" heatid="29008" />
                <RESULT resultid="5047" eventid="31" swimtime="00:01:12.43" lane="7" heatid="31002" />
                <RESULT resultid="5048" eventid="33" swimtime="00:01:46.18" lane="7" heatid="33003" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1081" birthdate="2014-01-01" gender="M" lastname="Polzin" firstname="Franz" license="451411">
              <RESULTS>
                <RESULT resultid="5049" eventid="22" swimtime="00:01:03.71" lane="5" heatid="22005" />
                <RESULT resultid="5050" eventid="26" swimtime="00:00:51.76" lane="6" heatid="26009" />
                <RESULT resultid="5051" eventid="30" swimtime="00:00:44.68" lane="1" heatid="30008" />
                <RESULT resultid="5052" eventid="32" swimtime="00:01:14.34" lane="1" heatid="32003" />
                <RESULT resultid="5053" eventid="34" swimtime="00:01:40.95" lane="7" heatid="34003" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1082" birthdate="2015-01-01" gender="F" lastname="Bindheim" firstname="Frieda" license="463477">
              <RESULTS>
                <RESULT resultid="5054" eventid="17" swimtime="00:01:16.34" lane="8" heatid="17003" />
                <RESULT resultid="5055" eventid="19" swimtime="00:01:12.39" lane="5" heatid="19002" />
                <RESULT resultid="5056" eventid="25" swimtime="00:01:00.81" lane="8" heatid="25004" />
                <RESULT resultid="5057" eventid="27" swimtime="00:01:23.61" lane="6" heatid="27001" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1083" birthdate="2009-01-01" gender="F" lastname="Rasmussen" firstname="Helen" license="398058">
              <RESULTS>
                <RESULT resultid="5058" eventid="5" swimtime="00:00:35.48" lane="2" heatid="5012" />
                <RESULT resultid="5059" eventid="10" swimtime="00:01:26.76" lane="3" heatid="10013" />
                <RESULT resultid="5060" eventid="12" swimtime="00:00:31.58" lane="7" heatid="12016" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1084" birthdate="2013-01-01" gender="M" lastname="Thiele" firstname="Henrik" license="451456">
              <RESULTS>
                <RESULT resultid="5061" eventid="4" swimtime="00:01:55.46" lane="8" heatid="4004" />
                <RESULT resultid="5062" eventid="11" swimtime="00:01:50.98" lane="6" heatid="11002" />
                <RESULT resultid="5063" eventid="13" swimtime="00:00:40.84" lane="6" heatid="13003" />
                <RESULT resultid="5064" eventid="20" swimtime="00:00:54.48" lane="1" heatid="20009" />
                <RESULT resultid="5065" eventid="26" swimtime="00:00:48.25" lane="5" heatid="26009" />
                <RESULT resultid="5066" eventid="28" swimtime="00:01:03.89" lane="7" heatid="28005" />
                <RESULT resultid="5067" eventid="34" swimtime="00:01:35.83" lane="3" heatid="34003" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1085" birthdate="2009-01-01" gender="M" lastname="Blazy" firstname="Janneck" license="421418">
              <RESULTS>
                <RESULT resultid="5068" eventid="20" swimtime="00:00:39.08" lane="6" heatid="20016" />
                <RESULT resultid="5069" eventid="24" swimtime="00:02:42.48" lane="5" heatid="24002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:15.81" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="5070" eventid="26" swimtime="00:00:36.26" lane="6" heatid="26020" />
                <RESULT resultid="5071" eventid="34" swimtime="00:01:10.78" lane="6" heatid="34011" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1086" birthdate="2015-01-01" gender="F" lastname="Hauschild" firstname="Julia" license="463480">
              <RESULTS>
                <RESULT resultid="5072" eventid="19" swimtime="00:01:03.26" lane="6" heatid="19004" />
                <RESULT resultid="5073" eventid="21" swimtime="00:01:36.16" lane="2" heatid="21002" />
                <RESULT resultid="5074" eventid="25" swimtime="00:01:00.85" lane="5" heatid="25003" />
                <RESULT resultid="5075" eventid="27" swimtime="00:01:23.07" lane="2" heatid="27001" />
                <RESULT resultid="5076" eventid="29" swimtime="00:00:56.43" lane="4" heatid="29003" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1087" birthdate="2014-01-01" gender="F" lastname="Brendler" firstname="Lena" license="451405">
              <RESULTS>
                <RESULT resultid="5077" eventid="21" swimtime="00:01:05.17" lane="5" heatid="21006" />
                <RESULT resultid="5078" eventid="25" swimtime="00:00:48.74" lane="8" heatid="25014" />
                <RESULT resultid="5079" eventid="29" swimtime="00:00:41.60" lane="2" heatid="29012" />
                <RESULT resultid="5080" eventid="31" swimtime="00:01:09.76" lane="1" heatid="31004" />
                <RESULT resultid="5081" eventid="33" swimtime="00:01:35.45" lane="1" heatid="33005" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1088" birthdate="2011-01-01" gender="F" lastname="Wilhelm" firstname="Linda" license="436850">
              <RESULTS>
                <RESULT resultid="5082" eventid="3" swimtime="00:01:45.19" lane="2" heatid="3006" />
                <RESULT resultid="5083" eventid="5" swimtime="00:00:42.65" lane="8" heatid="5008" />
                <RESULT resultid="5084" eventid="10" swimtime="00:01:30.94" lane="3" heatid="10010" />
                <RESULT resultid="5085" eventid="12" swimtime="00:00:35.28" lane="5" heatid="12009" />
                <RESULT resultid="5086" eventid="19" swimtime="00:00:47.27" lane="6" heatid="19017" />
                <RESULT resultid="5087" eventid="25" swimtime="00:00:41.63" lane="5" heatid="25025" />
                <RESULT resultid="5088" eventid="33" swimtime="00:01:20.62" lane="7" heatid="33011" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1089" birthdate="2015-01-01" gender="F" lastname="Heinitz" firstname="Linn" license="467472">
              <RESULTS>
                <RESULT resultid="5089" eventid="17" swimtime="00:01:26.01" lane="3" heatid="17007" />
                <RESULT resultid="5090" eventid="19" swimtime="00:01:00.53" lane="4" heatid="19010" />
                <RESULT resultid="5091" eventid="21" swimtime="00:01:11.61" lane="1" heatid="21006" />
                <RESULT resultid="5092" eventid="25" swimtime="00:00:55.98" lane="5" heatid="25008" />
                <RESULT resultid="5093" eventid="29" swimtime="00:00:47.09" lane="8" heatid="29010" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1090" birthdate="2013-01-01" gender="F" lastname="Sehr" firstname="Liska Amelia" license="444105">
              <RESULTS>
                <RESULT resultid="5094" eventid="3" swimtime="00:01:54.76" lane="2" heatid="3004" />
                <RESULT resultid="5095" eventid="12" swimtime="00:00:45.95" lane="2" heatid="12002" />
                <RESULT resultid="5096" eventid="19" swimtime="00:00:51.83" lane="6" heatid="19014" />
                <RESULT resultid="5097" eventid="25" swimtime="00:00:49.84" lane="3" heatid="25015" />
                <RESULT resultid="5098" eventid="27" swimtime="00:01:00.42" lane="5" heatid="27009" />
                <RESULT resultid="5099" eventid="31" swimtime="00:01:05.27" lane="8" heatid="31004" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1091" birthdate="2014-01-01" gender="F" lastname="Möbius" firstname="Lotte" license="451461">
              <RESULTS>
                <RESULT resultid="5100" eventid="17" swimtime="00:01:04.72" lane="2" heatid="17011" />
                <RESULT resultid="5101" eventid="19" swimtime="00:00:58.53" lane="8" heatid="19010" />
                <RESULT resultid="5102" eventid="25" swimtime="00:00:51.92" lane="4" heatid="25010" />
                <RESULT resultid="5103" eventid="29" swimtime="00:00:44.36" lane="5" heatid="29009" />
                <RESULT resultid="5104" eventid="31" swimtime="00:01:11.37" lane="7" heatid="31003" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1092" birthdate="2012-01-01" gender="F" lastname="Wandschneider" firstname="Marie" license="436844">
              <RESULTS>
                <RESULT resultid="5105" eventid="5" swimtime="00:00:48.93" lane="5" heatid="5003" />
                <RESULT resultid="5106" eventid="10" swimtime="00:01:43.33" lane="6" heatid="10005" />
                <RESULT resultid="5107" eventid="12" swimtime="00:00:43.30" lane="5" heatid="12004" />
                <RESULT resultid="5108" eventid="17" swimtime="00:01:00.73" lane="1" heatid="17012" />
                <RESULT resultid="5109" eventid="25" swimtime="00:00:46.78" lane="1" heatid="25020" />
                <RESULT resultid="5110" eventid="31" swimtime="00:00:59.99" lane="5" heatid="31005" />
                <RESULT resultid="5111" eventid="33" swimtime="00:01:27.96" lane="2" heatid="33007" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1093" birthdate="2014-01-01" gender="F" lastname="Huerta-Stiehl" firstname="Nelly Johanna" license="451404">
              <RESULTS>
                <RESULT resultid="5112" eventid="19" swimtime="00:00:52.61" lane="4" heatid="19015" />
                <RESULT resultid="5113" eventid="25" swimtime="00:00:55.32" lane="5" heatid="25009" />
                <RESULT resultid="5114" eventid="27" swimtime="00:01:03.25" lane="7" heatid="27006" />
                <RESULT resultid="5115" eventid="29" swimtime="00:00:47.33" lane="6" heatid="29007" />
                <RESULT resultid="5116" eventid="33" swimtime="00:01:47.91" lane="5" heatid="33002" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1094" birthdate="2015-01-01" gender="F" lastname="Dozsa-Nemeth" firstname="Odett" license="463478">
              <RESULTS>
                <RESULT resultid="5117" eventid="17" status="DNS" swimtime="00:00:00.00" lane="8" heatid="17009" />
                <RESULT resultid="5118" eventid="19" swimtime="00:01:00.80" lane="7" heatid="19007" />
                <RESULT resultid="5119" eventid="25" swimtime="00:00:51.94" lane="6" heatid="25015" />
                <RESULT resultid="5120" eventid="27" swimtime="00:01:15.91" lane="8" heatid="27005" />
                <RESULT resultid="5121" eventid="29" swimtime="00:00:46.57" lane="1" heatid="29010" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1095" birthdate="2015-01-01" gender="F" lastname="Naumann" firstname="Phyllis Maira" license="463481">
              <RESULTS>
                <RESULT resultid="5122" eventid="17" swimtime="00:01:17.80" lane="4" heatid="17002" />
                <RESULT resultid="5123" eventid="19" swimtime="00:01:09.86" lane="2" heatid="19003" />
                <RESULT resultid="5124" eventid="25" swimtime="00:01:05.42" lane="7" heatid="25003" />
                <RESULT resultid="5125" eventid="29" swimtime="00:00:59.35" lane="5" heatid="29003" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1096" birthdate="2015-01-01" gender="F" lastname="Otto" firstname="Pia" license="463476">
              <RESULTS>
                <RESULT resultid="5126" eventid="17" swimtime="00:01:00.20" lane="4" heatid="17010" />
                <RESULT resultid="5127" eventid="19" swimtime="00:00:57.56" lane="1" heatid="19014" />
                <RESULT resultid="5128" eventid="25" swimtime="00:00:48.07" lane="2" heatid="25020" />
                <RESULT resultid="5129" eventid="27" swimtime="00:01:08.94" lane="6" heatid="27006" />
                <RESULT resultid="5130" eventid="29" swimtime="00:00:43.00" lane="6" heatid="29012" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1097" birthdate="2007-01-01" gender="M" lastname="Maneck" firstname="Samuel" license="405759">
              <RESULTS>
                <RESULT resultid="5131" eventid="2" swimtime="00:02:35.14" lane="1" heatid="2008">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:09.79" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="5132" eventid="6" swimtime="00:00:27.53" lane="5" heatid="6011" />
                <RESULT resultid="5133" eventid="11" swimtime="00:01:11.23" lane="7" heatid="11012" />
                <RESULT resultid="5134" eventid="13" swimtime="00:00:26.57" lane="3" heatid="13018" />
                <RESULT resultid="5135" eventid="20" swimtime="00:00:35.33" lane="7" heatid="20022" />
                <RESULT resultid="5136" eventid="24" swimtime="00:02:15.50" lane="6" heatid="24009">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:05.41" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="5137" eventid="34" swimtime="00:00:59.04" lane="5" heatid="34015" />
                <RESULT resultid="5138" eventid="36" swimtime="00:01:07.31" lane="5" heatid="36003" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1098" birthdate="2013-01-01" gender="F" lastname="Voigt" firstname="Sophia" license="444104">
              <RESULTS>
                <RESULT resultid="5139" eventid="5" swimtime="00:00:51.21" lane="8" heatid="5003" />
                <RESULT resultid="5140" eventid="10" swimtime="00:01:29.14" lane="8" heatid="10011" />
                <RESULT resultid="5141" eventid="12" swimtime="00:00:35.69" lane="7" heatid="12010" />
                <RESULT resultid="5142" eventid="21" swimtime="00:00:51.01" lane="6" heatid="21014" />
                <RESULT resultid="5143" eventid="25" swimtime="00:00:41.69" lane="3" heatid="25023" />
                <RESULT resultid="5144" eventid="33" swimtime="00:01:19.36" lane="8" heatid="33013" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1099" birthdate="2011-01-01" gender="F" lastname="Harbich" firstname="Svea" license="422683">
              <RESULTS>
                <RESULT resultid="5145" eventid="3" swimtime="00:01:37.35" lane="8" heatid="3010" />
                <RESULT resultid="5146" eventid="10" swimtime="00:01:30.68" lane="5" heatid="10011" />
                <RESULT resultid="5147" eventid="12" swimtime="00:00:35.60" lane="8" heatid="12013" />
                <RESULT resultid="5148" eventid="19" swimtime="00:00:45.20" lane="5" heatid="19025" />
                <RESULT resultid="5149" eventid="25" swimtime="00:00:41.61" lane="2" heatid="25030" />
                <RESULT resultid="5150" eventid="33" swimtime="00:01:19.45" lane="3" heatid="33014" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1100" birthdate="2011-01-01" gender="F" lastname="Duckstein" firstname="Tanja" license="422686">
              <RESULTS>
                <RESULT resultid="5151" eventid="23" swimtime="00:02:39.66" lane="4" heatid="23009">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:18.14" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="5152" eventid="33" swimtime="00:01:13.73" lane="4" heatid="33016" />
                <RESULT resultid="5153" eventid="35" swimtime="00:01:29.55" lane="3" heatid="35003" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1102" birthdate="2013-01-01" gender="F" lastname="Voigt" firstname="Victoria" license="444805">
              <RESULTS>
                <RESULT resultid="5161" eventid="3" swimtime="00:01:58.24" lane="4" heatid="3003" />
                <RESULT resultid="5162" eventid="12" swimtime="00:00:45.61" lane="1" heatid="12006" />
                <RESULT resultid="5163" eventid="17" status="DNS" swimtime="00:00:00.00" lane="2" heatid="17012" />
                <RESULT resultid="5164" eventid="19" status="DNS" swimtime="00:00:00.00" lane="6" heatid="19012" />
                <RESULT resultid="5165" eventid="27" status="DNS" swimtime="00:00:00.00" lane="8" heatid="27010" />
                <RESULT resultid="5166" eventid="33" status="DNS" swimtime="00:00:00.00" lane="3" heatid="33006" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1103" birthdate="2012-01-01" gender="M" lastname="Stäudte" firstname="Vincent" license="436853">
              <RESULTS>
                <RESULT resultid="5167" eventid="4" swimtime="00:01:37.76" lane="3" heatid="4008" />
                <RESULT resultid="5168" eventid="6" swimtime="00:00:36.26" lane="2" heatid="6008" />
                <RESULT resultid="5169" eventid="11" swimtime="00:01:19.30" lane="5" heatid="11011" />
                <RESULT resultid="5170" eventid="13" swimtime="00:00:32.50" lane="7" heatid="13013" />
                <RESULT resultid="5171" eventid="24" swimtime="00:02:32.27" lane="7" heatid="24008">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:13.46" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="5172" eventid="26" swimtime="00:00:35.49" lane="2" heatid="26022" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1104" birthdate="2013-01-01" gender="M" lastname="Geleschus" firstname="Yannick" license="449831">
              <RESULTS>
                <RESULT resultid="5173" eventid="22" swimtime="00:00:55.22" lane="2" heatid="22010" />
                <RESULT resultid="5174" eventid="24" swimtime="00:03:12.16" lane="8" heatid="24003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:34.34" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="5175" eventid="32" swimtime="00:00:59.42" lane="2" heatid="32004" />
                <RESULT resultid="5176" eventid="34" swimtime="00:01:30.43" lane="2" heatid="34005" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1105" birthdate="2012-01-01" gender="F" lastname="Kobsik" firstname="Zoe" license="449834">
              <RESULTS>
                <RESULT resultid="5177" eventid="5" swimtime="00:00:39.33" lane="7" heatid="5007" />
                <RESULT resultid="5178" eventid="10" swimtime="00:01:38.33" lane="7" heatid="10009" />
                <RESULT resultid="5179" eventid="12" swimtime="00:00:33.97" lane="8" heatid="12011" />
                <RESULT resultid="5180" eventid="17" swimtime="00:00:54.14" lane="6" heatid="17015" />
                <RESULT resultid="5181" eventid="21" swimtime="00:00:50.79" lane="4" heatid="21013" />
                <RESULT resultid="5182" eventid="33" swimtime="00:01:15.87" lane="4" heatid="33013" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="SV 1990 Zschopau" nation="GER" region="12" code="3382">
          <ATHLETES>
            <ATHLETE athleteid="992" birthdate="2013-01-01" gender="F" lastname="Keller" firstname="Emma" license="460563">
              <RESULTS>
                <RESULT resultid="4613" eventid="3" swimtime="00:01:58.23" lane="3" heatid="3003" />
                <RESULT resultid="4614" eventid="5" swimtime="00:00:46.99" lane="5" heatid="5004" />
                <RESULT resultid="4615" eventid="10" status="DNS" swimtime="00:00:00.00" lane="5" heatid="10001" />
                <RESULT resultid="4616" eventid="12" swimtime="00:00:40.11" lane="8" heatid="12006" />
                <RESULT resultid="4617" eventid="19" swimtime="00:00:54.44" lane="3" heatid="19014" />
                <RESULT resultid="4618" eventid="21" swimtime="00:00:57.06" lane="7" heatid="21013" />
                <RESULT resultid="4619" eventid="27" swimtime="00:01:11.60" lane="3" heatid="27001" />
                <RESULT resultid="4620" eventid="31" swimtime="00:01:00.53" lane="4" heatid="31005" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="993" birthdate="2007-01-01" gender="F" lastname="Tanneberger" firstname="Fiona" license="430278">
              <RESULTS>
                <RESULT resultid="4621" eventid="3" swimtime="00:01:30.52" lane="7" heatid="3011" />
                <RESULT resultid="4622" eventid="10" swimtime="00:01:25.11" lane="4" heatid="10010" />
                <RESULT resultid="4623" eventid="12" swimtime="00:00:31.17" lane="7" heatid="12015" />
                <RESULT resultid="4624" eventid="14" swimtime="00:03:22.20" lane="4" heatid="14006">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:38.29" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="994" birthdate="2010-01-01" gender="M" lastname="Zingler" firstname="Gustav Albert" license="409207">
              <RESULTS>
                <RESULT resultid="4625" eventid="4" swimtime="00:01:24.05" lane="2" heatid="4011" />
                <RESULT resultid="4626" eventid="6" swimtime="00:00:31.94" lane="8" heatid="6010" />
                <RESULT resultid="4627" eventid="13" swimtime="00:00:29.54" lane="5" heatid="13016" />
                <RESULT resultid="4628" eventid="15" swimtime="00:03:11.90" lane="7" heatid="15007">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:32.17" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="4629" eventid="20" swimtime="00:00:36.39" lane="3" heatid="20022" />
                <RESULT resultid="4630" eventid="24" swimtime="00:02:34.04" lane="4" heatid="24008">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:11.60" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="4631" eventid="34" swimtime="00:01:06.97" lane="2" heatid="34014" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="995" birthdate="2013-01-01" gender="F" lastname="Decker" firstname="Helene" license="464574">
              <RESULTS>
                <RESULT resultid="4632" eventid="3" swimtime="00:02:01.12" lane="6" heatid="3003" />
                <RESULT resultid="4633" eventid="10" swimtime="00:01:50.10" lane="4" heatid="10002" />
                <RESULT resultid="4634" eventid="12" swimtime="00:00:43.37" lane="5" heatid="12003" />
                <RESULT resultid="4635" eventid="17" swimtime="00:01:07.92" lane="1" heatid="17006" />
                <RESULT resultid="4636" eventid="19" swimtime="00:00:56.91" lane="6" heatid="19013" />
                <RESULT resultid="4637" eventid="25" swimtime="00:00:50.08" lane="5" heatid="25017" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="996" birthdate="2011-01-01" gender="M" lastname="Schmieder" firstname="Julian Magnus" license="394210">
              <RESULTS>
                <RESULT resultid="4638" eventid="4" swimtime="00:01:59.89" lane="6" heatid="4003" />
                <RESULT resultid="4639" eventid="11" swimtime="00:01:41.08" lane="1" heatid="11005" />
                <RESULT resultid="4640" eventid="13" swimtime="00:00:39.57" lane="6" heatid="13004" />
                <RESULT resultid="4641" eventid="20" swimtime="00:00:54.78" lane="4" heatid="20008" />
                <RESULT resultid="4642" eventid="26" swimtime="00:00:45.68" lane="3" heatid="26014" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="997" birthdate="2014-01-01" gender="F" lastname="Meusel" firstname="Lotta Chayenne" license="474377">
              <RESULTS>
                <RESULT resultid="4643" eventid="17" swimtime="00:01:22.19" lane="7" heatid="17001" />
                <RESULT resultid="4644" eventid="19" status="DSQ" swimtime="00:01:06.25" lane="4" heatid="19003" comment="Start vor dem Startsignal." />
                <RESULT resultid="4645" eventid="25" swimtime="00:01:06.12" lane="1" heatid="25003" />
                <RESULT resultid="4646" eventid="29" swimtime="00:01:07.68" lane="6" heatid="29002" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="998" birthdate="2007-01-01" gender="F" lastname="Zingler" firstname="Lotte Pauline" license="365814">
              <RESULTS>
                <RESULT resultid="4647" eventid="1" swimtime="00:02:58.76" lane="3" heatid="1004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:21.19" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="4648" eventid="5" swimtime="00:00:35.46" lane="1" heatid="5012" />
                <RESULT resultid="4649" eventid="10" swimtime="00:01:22.65" lane="5" heatid="10015" />
                <RESULT resultid="4650" eventid="12" swimtime="00:00:32.18" lane="5" heatid="12016" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="999" birthdate="2007-01-01" gender="F" lastname="Guba" firstname="Mailin" license="393192">
              <RESULTS>
                <RESULT resultid="4651" eventid="19" swimtime="00:00:47.20" lane="6" heatid="19023" />
                <RESULT resultid="4652" eventid="23" swimtime="00:02:55.12" lane="2" heatid="23004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:20.76" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="4653" eventid="33" swimtime="00:01:16.45" lane="5" heatid="33015" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1000" birthdate="2014-01-01" gender="M" lastname="Reuter" firstname="Nils" license="464573">
              <RESULTS>
                <RESULT resultid="4654" eventid="20" swimtime="00:00:56.61" lane="5" heatid="20005" />
                <RESULT resultid="4655" eventid="26" swimtime="00:00:57.18" lane="6" heatid="26011" />
                <RESULT resultid="4656" eventid="28" swimtime="00:01:13.71" lane="6" heatid="28001" />
                <RESULT resultid="4657" eventid="30" swimtime="00:00:44.11" lane="8" heatid="30007" />
                <RESULT resultid="4658" eventid="32" swimtime="00:01:13.15" lane="7" heatid="32002" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1001" birthdate="2008-01-01" gender="M" lastname="Meusel" firstname="Noah Joel" license="393191">
              <RESULTS>
                <RESULT resultid="4659" eventid="4" swimtime="00:01:31.99" lane="5" heatid="4009" />
                <RESULT resultid="4660" eventid="6" swimtime="00:00:31.77" lane="3" heatid="6010" />
                <RESULT resultid="4661" eventid="13" swimtime="00:00:29.78" lane="6" heatid="13016" />
                <RESULT resultid="4662" eventid="20" swimtime="00:00:39.09" lane="2" heatid="20021" />
                <RESULT resultid="4663" eventid="24" swimtime="00:02:34.54" lane="4" heatid="24007">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:13.29" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="4664" eventid="34" swimtime="00:01:05.35" lane="6" heatid="34014" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="SV Automation e.V." nation="GER" region="12" code="6435">
          <ATHLETES>
            <ATHLETE athleteid="436" birthdate="2012-01-01" gender="M" lastname="Birgel" firstname="Mick" license="407310">
              <RESULTS>
                <RESULT resultid="2109" eventid="2" swimtime="00:02:54.22" lane="1" heatid="2006">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:22.66" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="2108" eventid="6" swimtime="00:00:35.32" lane="8" heatid="6008" />
                <RESULT resultid="2107" eventid="11" swimtime="00:01:19.85" lane="4" heatid="11009" />
                <RESULT resultid="2106" eventid="13" swimtime="00:00:32.21" lane="7" heatid="13012" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="437" birthdate="2012-01-01" gender="M" lastname="Sauerteig" firstname="Johann" license="434534">
              <RESULTS>
                <RESULT resultid="2113" eventid="4" status="DSQ" swimtime="00:01:47.48" lane="8" heatid="4005" comment="Start vor dem Startsignal." />
                <RESULT resultid="2112" eventid="6" swimtime="00:00:57.79" lane="5" heatid="6002" />
                <RESULT resultid="2111" eventid="11" swimtime="00:01:52.76" lane="1" heatid="11003" />
                <RESULT resultid="2110" eventid="13" swimtime="00:00:41.07" lane="2" heatid="13003" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="438" birthdate="2012-01-01" gender="F" lastname="Janz" firstname="Joanne Savannah" license="424375">
              <RESULTS>
                <RESULT resultid="2116" eventid="3" swimtime="00:01:45.01" lane="7" heatid="3005" />
                <RESULT resultid="2115" eventid="10" swimtime="00:01:35.00" lane="3" heatid="10005" />
                <RESULT resultid="2114" eventid="12" swimtime="00:00:38.49" lane="7" heatid="12008" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="439" birthdate="2012-01-01" gender="M" lastname="Szabo" firstname="Janos" license="440685">
              <RESULTS>
                <RESULT resultid="2120" eventid="4" swimtime="00:01:47.14" lane="5" heatid="4004" />
                <RESULT resultid="2119" eventid="6" swimtime="00:00:44.26" lane="4" heatid="6002" />
                <RESULT resultid="2118" eventid="11" swimtime="00:01:27.59" lane="1" heatid="11006" />
                <RESULT resultid="2117" eventid="13" swimtime="00:00:36.41" lane="8" heatid="13007" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="440" birthdate="2013-01-01" gender="F" lastname="Münchhof" firstname="Ina" license="445227">
              <RESULTS>
                <RESULT resultid="2123" eventid="5" swimtime="00:00:44.08" lane="8" heatid="5007" />
                <RESULT resultid="2122" eventid="10" swimtime="00:01:36.35" lane="4" heatid="10005" />
                <RESULT resultid="2121" eventid="12" swimtime="00:00:37.81" lane="6" heatid="12004" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="441" birthdate="2012-01-01" gender="F" lastname="Wießner" firstname="Emilia" license="434536">
              <RESULTS>
                <RESULT resultid="2127" eventid="1" swimtime="00:03:08.60" lane="8" heatid="1004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:29.24" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="2126" eventid="3" swimtime="00:01:40.45" lane="6" heatid="3007" />
                <RESULT resultid="2125" eventid="10" swimtime="00:01:27.04" lane="4" heatid="10007" />
                <RESULT resultid="2124" eventid="12" swimtime="00:00:34.47" lane="1" heatid="12013" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="442" birthdate="2013-01-01" gender="M" lastname="Hottas" firstname="Casper" license="440671">
              <RESULTS>
                <RESULT resultid="2131" eventid="18" swimtime="00:01:02.13" lane="7" heatid="18008" />
                <RESULT resultid="2130" eventid="24" swimtime="00:03:35.67" lane="6" heatid="24002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:44.75" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="2129" eventid="32" swimtime="00:00:58.49" lane="4" heatid="32004" />
                <RESULT resultid="2128" eventid="36" swimtime="00:01:50.24" lane="4" heatid="36001" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="443" birthdate="2012-01-01" gender="M" lastname="Zens" firstname="Caspar Valentin" license="444869">
              <RESULTS>
                <RESULT resultid="2135" eventid="22" swimtime="00:00:48.96" lane="2" heatid="22011" />
                <RESULT resultid="2134" eventid="24" swimtime="00:02:47.59" lane="7" heatid="24007">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:21.60" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="2133" eventid="32" swimtime="00:00:53.48" lane="2" heatid="32005" />
                <RESULT resultid="2132" eventid="36" swimtime="00:01:29.96" lane="2" heatid="36002" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="444" birthdate="2011-01-01" gender="F" lastname="Dyka" firstname="Arina" license="456586">
              <RESULTS>
                <RESULT resultid="2143" eventid="1" swimtime="00:02:50.03" lane="8" heatid="1007">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:21.25" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="2142" eventid="5" swimtime="00:00:34.81" lane="5" heatid="5011" />
                <RESULT resultid="2141" eventid="8" swimtime="00:03:06.27" lane="3" heatid="8001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:24.87" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="2140" eventid="12" swimtime="00:00:32.29" lane="1" heatid="12016" />
                <RESULT resultid="2139" eventid="19" swimtime="00:00:40.47" lane="7" heatid="19026" />
                <RESULT resultid="2138" eventid="25" swimtime="00:00:38.49" lane="8" heatid="25029" />
                <RESULT resultid="2137" eventid="33" swimtime="00:01:09.36" lane="2" heatid="33017" />
                <RESULT resultid="2136" eventid="37" swimtime="00:02:54.30" lane="7" heatid="37005">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:26.13" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="SV Dresden-Nord" nation="GER" region="12" code="3386">
          <ATHLETES>
            <ATHLETE athleteid="87" birthdate="2013-01-01" gender="F" lastname="Schwendler" firstname="Alexandra" license="449958">
              <RESULTS>
                <RESULT resultid="470" eventid="3" swimtime="00:01:53.76" lane="8" heatid="3003" />
                <RESULT resultid="471" eventid="10" status="DSQ" swimtime="00:01:42.40" lane="2" heatid="10004" comment="Nach verlassen der Rückenlage Wende nicht unverzüglich eingeleitet." />
                <RESULT resultid="472" eventid="12" swimtime="00:00:37.77" lane="2" heatid="12006" />
                <RESULT resultid="473" eventid="17" swimtime="00:00:52.33" lane="6" heatid="17016" />
                <RESULT resultid="474" eventid="25" swimtime="00:00:45.57" lane="6" heatid="25022" />
                <RESULT resultid="475" eventid="31" swimtime="00:00:59.30" lane="5" heatid="31002" />
                <RESULT resultid="476" eventid="33" swimtime="00:01:27.94" lane="4" heatid="33005" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="88" birthdate="2014-01-01" gender="M" lastname="Olbrich" firstname="Max" license="474578">
              <RESULTS>
                <RESULT resultid="477" eventid="20" swimtime="00:00:56.50" lane="1" heatid="20008" />
                <RESULT resultid="478" eventid="22" swimtime="00:01:03.34" lane="4" heatid="22002" />
                <RESULT resultid="479" eventid="26" swimtime="00:00:55.80" lane="7" heatid="26010" />
                <RESULT resultid="480" eventid="28" swimtime="00:01:05.21" lane="2" heatid="28002" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="SV Fortschritt Pirna" nation="GER" region="12" code="3387">
          <ATHLETES>
            <ATHLETE athleteid="878" birthdate="2012-01-01" gender="M" lastname="Adler" firstname="Bendix" license="448850">
              <RESULTS>
                <RESULT resultid="4111" eventid="11" swimtime="00:01:24.95" lane="3" heatid="11004" />
                <RESULT resultid="4112" eventid="13" swimtime="00:00:32.25" lane="5" heatid="13011" />
                <RESULT resultid="4113" eventid="15" swimtime="00:03:14.78" lane="4" heatid="15005">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:32.54" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="4114" eventid="24" swimtime="00:02:42.05" lane="6" heatid="24007">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:17.71" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="879" birthdate="2014-01-01" gender="M" lastname="Tanner" firstname="German" license="457699">
              <RESULTS>
                <RESULT resultid="4115" eventid="18" swimtime="00:01:06.68" lane="3" heatid="18004" />
                <RESULT resultid="4116" eventid="20" swimtime="00:01:02.77" lane="1" heatid="20004" />
                <RESULT resultid="4117" eventid="22" swimtime="00:01:08.12" lane="1" heatid="22004" />
                <RESULT resultid="4118" eventid="26" status="DSQ" swimtime="00:00:53.30" lane="3" heatid="26005" comment="Start vor dem Startsignal." />
                <RESULT resultid="4119" eventid="30" swimtime="00:00:46.21" lane="6" heatid="30004" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="880" birthdate="2014-01-01" gender="F" lastname="Hein" firstname="Helen Ronja" license="448835">
              <RESULTS>
                <RESULT resultid="4120" eventid="19" swimtime="00:00:56.37" lane="8" heatid="19009" />
                <RESULT resultid="4121" eventid="21" swimtime="00:00:53.58" lane="8" heatid="21014" />
                <RESULT resultid="4122" eventid="29" swimtime="00:00:40.19" lane="5" heatid="29008" />
                <RESULT resultid="4123" eventid="31" swimtime="00:01:00.13" lane="2" heatid="31005" />
                <RESULT resultid="4124" eventid="33" swimtime="00:01:39.74" lane="4" heatid="33004" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="881" birthdate="2013-01-01" gender="F" lastname="Kirsch" firstname="Hermine" license="452328">
              <RESULTS>
                <RESULT resultid="4125" eventid="3" swimtime="00:02:11.81" lane="5" heatid="3001" />
                <RESULT resultid="4126" eventid="10" swimtime="00:01:58.68" lane="4" heatid="10001" />
                <RESULT resultid="4127" eventid="12" swimtime="00:00:44.97" lane="4" heatid="12001" />
                <RESULT resultid="4128" eventid="19" swimtime="00:01:01.15" lane="5" heatid="19004" />
                <RESULT resultid="4129" eventid="21" swimtime="00:01:11.13" lane="7" heatid="21004" />
                <RESULT resultid="4130" eventid="27" swimtime="00:01:11.39" lane="8" heatid="27004" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="882" birthdate="2011-01-01" gender="F" lastname="Schoss" firstname="Johanna" license="437047">
              <RESULTS>
                <RESULT resultid="4131" eventid="3" swimtime="00:01:55.12" lane="4" heatid="3002" />
                <RESULT resultid="4132" eventid="10" status="DNS" swimtime="00:00:00.00" lane="8" heatid="10003" />
                <RESULT resultid="4133" eventid="12" swimtime="00:00:38.40" lane="5" heatid="12006" />
                <RESULT resultid="4134" eventid="19" status="DNS" swimtime="00:00:00.00" lane="6" heatid="19015" />
                <RESULT resultid="4135" eventid="25" status="DNS" swimtime="00:00:00.00" lane="5" heatid="25020" />
                <RESULT resultid="4136" eventid="33" status="DNS" swimtime="00:00:00.00" lane="8" heatid="33004" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="883" birthdate="2014-01-01" gender="F" lastname="Wittka" firstname="Johanna" license="457673">
              <RESULTS>
                <RESULT resultid="4137" eventid="17" swimtime="00:01:08.56" lane="5" heatid="17001" />
                <RESULT resultid="4138" eventid="19" swimtime="00:01:02.59" lane="1" heatid="19005" />
                <RESULT resultid="4139" eventid="21" swimtime="00:00:59.81" lane="3" heatid="21005" />
                <RESULT resultid="4140" eventid="25" swimtime="00:00:53.38" lane="2" heatid="25009" />
                <RESULT resultid="4141" eventid="29" swimtime="00:00:45.91" lane="8" heatid="29006" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="884" birthdate="2014-01-01" gender="M" lastname="Schoss" firstname="Karl" license="448834">
              <RESULTS>
                <RESULT resultid="4142" eventid="18" swimtime="00:01:05.29" lane="3" heatid="18008" />
                <RESULT resultid="4143" eventid="22" swimtime="00:00:54.02" lane="7" heatid="22010" />
                <RESULT resultid="4144" eventid="30" swimtime="00:00:41.65" lane="3" heatid="30006" />
                <RESULT resultid="4145" eventid="32" swimtime="00:01:01.00" lane="2" heatid="32003" />
                <RESULT resultid="4146" eventid="34" swimtime="00:01:52.89" lane="4" heatid="34001" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="885" birthdate="2014-01-01" gender="F" lastname="Kaiser" firstname="Laura" license="460046">
              <RESULTS>
                <RESULT resultid="4147" eventid="17" status="DSQ" swimtime="00:01:15.83" lane="7" heatid="17004" comment="Start vor dem Startsignal." />
                <RESULT resultid="4148" eventid="19" swimtime="00:01:01.72" lane="7" heatid="19006" />
                <RESULT resultid="4149" eventid="25" status="DSQ" swimtime="00:00:55.15" lane="4" heatid="25009" comment="Start vor dem Startsignal." />
                <RESULT resultid="4150" eventid="27" swimtime="00:01:11.80" lane="4" heatid="27004" />
                <RESULT resultid="4151" eventid="29" swimtime="00:00:49.51" lane="1" heatid="29004" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="886" birthdate="2015-01-01" gender="F" lastname="Hofmann" firstname="Lucy" license="475224">
              <RESULTS>
                <RESULT resultid="4152" eventid="17" status="DSQ" swimtime="00:00:57.08" lane="1" heatid="17002" comment="Rücken Gesamtbewegung geschwommen." />
                <RESULT resultid="4153" eventid="19" status="DSQ" swimtime="00:01:04.82" lane="7" heatid="19003" comment="Der Zielanschlag erfolgte nur mit einer Hand." />
                <RESULT resultid="4154" eventid="21" swimtime="00:01:08.09" lane="5" heatid="21003" />
                <RESULT resultid="4155" eventid="25" swimtime="00:00:56.31" lane="2" heatid="25002" />
                <RESULT resultid="4156" eventid="29" swimtime="00:00:51.82" lane="8" heatid="29003" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="887" birthdate="2013-01-01" gender="F" lastname="Lindenmüller" firstname="Mara" license="448838">
              <RESULTS>
                <RESULT resultid="4157" eventid="3" swimtime="00:02:10.55" lane="3" heatid="3001" />
                <RESULT resultid="4158" eventid="10" swimtime="00:01:52.74" lane="7" heatid="10002" />
                <RESULT resultid="4159" eventid="12" swimtime="00:00:46.19" lane="3" heatid="12002" />
                <RESULT resultid="4160" eventid="19" swimtime="00:01:01.43" lane="1" heatid="19004" />
                <RESULT resultid="4161" eventid="21" swimtime="00:01:18.56" lane="6" heatid="21002" />
                <RESULT resultid="4162" eventid="27" swimtime="00:01:12.12" lane="7" heatid="27004" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="888" birthdate="2015-01-01" gender="M" lastname="Wittka" firstname="Oskar" license="475221">
              <RESULTS>
                <RESULT resultid="4163" eventid="18" swimtime="00:01:10.35" lane="5" heatid="18002" />
                <RESULT resultid="4164" eventid="22" swimtime="00:01:01.99" lane="7" heatid="22005" />
                <RESULT resultid="4165" eventid="26" swimtime="00:01:00.09" lane="5" heatid="26001" />
                <RESULT resultid="4166" eventid="30" status="DNS" swimtime="00:00:00.00" lane="1" heatid="30001" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="889" birthdate="2012-01-01" gender="M" lastname="Tobias" firstname="René Franz" license="448831">
              <RESULTS>
                <RESULT resultid="4167" eventid="4" swimtime="00:02:09.81" lane="5" heatid="4001" />
                <RESULT resultid="4168" eventid="11" swimtime="00:01:56.56" lane="7" heatid="11002" />
                <RESULT resultid="4169" eventid="13" swimtime="00:00:43.31" lane="3" heatid="13002" />
                <RESULT resultid="4170" eventid="20" swimtime="00:00:59.33" lane="6" heatid="20001" />
                <RESULT resultid="4171" eventid="22" swimtime="00:01:00.18" lane="6" heatid="22006" />
                <RESULT resultid="4172" eventid="28" status="DSQ" swimtime="00:01:06.18" lane="4" heatid="28002" comment="Das Brett wurde beim Anschlag vorn nicht umfasst." />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="890" birthdate="2013-01-01" gender="M" lastname="Gruhl" firstname="Theodor" license="445434">
              <RESULTS>
                <RESULT resultid="4173" eventid="2" swimtime="00:03:55.69" lane="4" heatid="2001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:48.91" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="4174" eventid="6" swimtime="00:00:44.69" lane="1" heatid="6002" />
                <RESULT resultid="4175" eventid="11" swimtime="00:01:44.14" lane="5" heatid="11001" />
                <RESULT resultid="4176" eventid="13" swimtime="00:00:37.86" lane="7" heatid="13004" />
                <RESULT resultid="4177" eventid="22" status="DSQ" swimtime="00:00:54.75" lane="8" heatid="22008" comment="Das Brett wurde beim Zielanschlag nicht umfasst." />
                <RESULT resultid="4178" eventid="26" swimtime="00:00:44.23" lane="7" heatid="26009" />
                <RESULT resultid="4179" eventid="34" swimtime="00:01:25.51" lane="7" heatid="34005" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="SV Handwerk Leipzig e.V." nation="GER" region="12" code="3390">
          <ATHLETES>
            <ATHLETE athleteid="892" birthdate="2015-01-01" gender="M" lastname="Gräfe" firstname="Adrian" license="467425">
              <RESULTS>
                <RESULT resultid="4184" eventid="18" swimtime="00:01:01.54" lane="6" heatid="18010" />
                <RESULT resultid="4185" eventid="22" swimtime="00:00:59.03" lane="7" heatid="22008" />
                <RESULT resultid="4186" eventid="26" swimtime="00:00:51.36" lane="4" heatid="26007" />
                <RESULT resultid="4187" eventid="30" swimtime="00:00:57.64" lane="5" heatid="30002" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="893" birthdate="2014-01-01" gender="M" lastname="Drechsel" firstname="Ben" license="449520">
              <RESULTS>
                <RESULT resultid="4188" eventid="18" swimtime="00:01:11.23" lane="1" heatid="18008" />
                <RESULT resultid="4189" eventid="20" swimtime="00:00:52.76" lane="5" heatid="20009" />
                <RESULT resultid="4190" eventid="22" swimtime="00:01:04.77" lane="1" heatid="22007" />
                <RESULT resultid="4191" eventid="28" swimtime="00:01:01.49" lane="3" heatid="28006" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="894" birthdate="2014-01-01" gender="M" lastname="Brückner" firstname="Carl" license="454910">
              <RESULTS>
                <RESULT resultid="4192" eventid="20" swimtime="00:00:54.23" lane="6" heatid="20007" />
                <RESULT resultid="4193" eventid="26" swimtime="00:00:45.64" lane="1" heatid="26012" />
                <RESULT resultid="4194" eventid="30" swimtime="00:00:41.05" lane="5" heatid="30007" />
                <RESULT resultid="4195" eventid="32" swimtime="00:01:00.15" lane="7" heatid="32004" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="895" birthdate="2014-01-01" gender="M" lastname="Suhayda" firstname="Ferdinand" license="449628">
              <RESULTS>
                <RESULT resultid="4196" eventid="20" swimtime="00:00:55.98" lane="2" heatid="20007" />
                <RESULT resultid="4197" eventid="22" swimtime="00:01:01.79" lane="5" heatid="22006" />
                <RESULT resultid="4198" eventid="26" swimtime="00:00:49.63" lane="1" heatid="26007" />
                <RESULT resultid="4199" eventid="28" swimtime="00:01:04.82" lane="3" heatid="28005" />
                <RESULT resultid="4200" eventid="30" swimtime="00:00:43.08" lane="4" heatid="30006" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="896" birthdate="2015-01-01" gender="F" lastname="Thomas" firstname="Hannah" license="460028">
              <RESULTS>
                <RESULT resultid="4201" eventid="17" swimtime="00:01:00.66" lane="5" heatid="17014" />
                <RESULT resultid="4202" eventid="21" swimtime="00:00:53.53" lane="3" heatid="21012" />
                <RESULT resultid="4203" eventid="25" swimtime="00:00:52.51" lane="1" heatid="25014" />
                <RESULT resultid="4204" eventid="29" swimtime="00:00:59.80" lane="5" heatid="29005" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="897" birthdate="2014-01-01" gender="M" lastname="Noack" firstname="Jakob" license="449525">
              <RESULTS>
                <RESULT resultid="4205" eventid="18" swimtime="00:00:56.01" lane="7" heatid="18011" />
                <RESULT resultid="4206" eventid="22" swimtime="00:00:56.31" lane="3" heatid="22009" />
                <RESULT resultid="4207" eventid="26" swimtime="00:00:48.05" lane="4" heatid="26010" />
                <RESULT resultid="4208" eventid="30" swimtime="00:00:46.98" lane="2" heatid="30005" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="898" birthdate="2014-01-01" gender="M" lastname="Engel" firstname="Johann" license="444263">
              <RESULTS>
                <RESULT resultid="4209" eventid="18" swimtime="00:01:19.21" lane="7" heatid="18002" />
                <RESULT resultid="4210" eventid="20" swimtime="00:00:49.00" lane="1" heatid="20012" />
                <RESULT resultid="4211" eventid="28" swimtime="00:00:57.56" lane="5" heatid="28007" />
                <RESULT resultid="4212" eventid="30" swimtime="00:00:48.78" lane="5" heatid="30005" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="899" birthdate="2014-01-01" gender="F" lastname="Schönwiesner" firstname="Jozefien" license="463049">
              <RESULTS>
                <RESULT resultid="4213" eventid="17" status="DNS" swimtime="00:00:00.00" lane="7" heatid="17012" />
                <RESULT resultid="4214" eventid="19" status="DNS" swimtime="00:00:00.00" lane="4" heatid="19002" />
                <RESULT resultid="4215" eventid="21" status="DNS" swimtime="00:00:00.00" lane="7" heatid="21006" />
                <RESULT resultid="4216" eventid="25" status="DNS" swimtime="00:00:00.00" lane="4" heatid="25013" />
                <RESULT resultid="4217" eventid="31" status="DNS" swimtime="00:00:00.00" lane="1" heatid="31002" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="900" birthdate="2015-01-01" gender="F" lastname="Leclerque" firstname="Judith" license="467426">
              <RESULTS>
                <RESULT resultid="4218" eventid="17" swimtime="00:01:07.80" lane="3" heatid="17005" />
                <RESULT resultid="4219" eventid="21" swimtime="00:01:05.49" lane="2" heatid="21006" />
                <RESULT resultid="4220" eventid="25" swimtime="00:00:57.18" lane="7" heatid="25005" />
                <RESULT resultid="4221" eventid="29" swimtime="00:00:58.67" lane="3" heatid="29002" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="901" birthdate="2015-01-01" gender="F" lastname="Herrmann Torres" firstname="Mia Hilde" license="467423">
              <RESULTS>
                <RESULT resultid="4222" eventid="17" swimtime="00:00:57.42" lane="8" heatid="17014" />
                <RESULT resultid="4223" eventid="21" swimtime="00:01:04.35" lane="7" heatid="21008" />
                <RESULT resultid="4224" eventid="25" swimtime="00:00:53.05" lane="8" heatid="25010" />
                <RESULT resultid="4225" eventid="29" swimtime="00:00:50.41" lane="2" heatid="29005" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="902" birthdate="2015-01-01" gender="F" lastname="Pinkau" firstname="Nadja" license="467427">
              <RESULTS>
                <RESULT resultid="4226" eventid="17" swimtime="00:01:03.99" lane="7" heatid="17011" />
                <RESULT resultid="4227" eventid="21" swimtime="00:01:02.26" lane="8" heatid="21008" />
                <RESULT resultid="4228" eventid="25" status="DSQ" swimtime="00:00:57.00" lane="6" heatid="25007" comment="Der Anschlag erfolgte nicht in Rückenlage." />
                <RESULT resultid="4229" eventid="27" swimtime="00:01:13.08" lane="1" heatid="27004" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="903" birthdate="2014-01-01" gender="M" lastname="Manitz" firstname="Paul Werner" license="457512">
              <RESULTS>
                <RESULT resultid="4230" eventid="18" swimtime="00:00:55.92" lane="4" heatid="18010" />
                <RESULT resultid="4231" eventid="26" swimtime="00:00:43.81" lane="5" heatid="26014" />
                <RESULT resultid="4232" eventid="30" swimtime="00:00:42.26" lane="2" heatid="30007" />
                <RESULT resultid="4233" eventid="32" swimtime="00:01:03.94" lane="5" heatid="32002" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="SV Lok Görlitz e.V." nation="GER" region="12" code="3337">
          <ATHLETES>
            <ATHLETE athleteid="1122" birthdate="2010-01-01" gender="F" lastname="Urban" firstname="Alisa Marie" license="415152">
              <RESULTS>
                <RESULT resultid="5255" eventid="3" swimtime="00:01:33.42" lane="2" heatid="3009" />
                <RESULT resultid="5256" eventid="12" swimtime="00:00:32.12" lane="4" heatid="12014" />
                <RESULT resultid="5257" eventid="14" swimtime="00:03:28.36" lane="7" heatid="14005">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:40.07" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1123" birthdate="2013-01-01" gender="M" lastname="Vogt" firstname="Aurelius" license="445775">
              <RESULTS>
                <RESULT resultid="5258" eventid="2" swimtime="00:03:31.69" lane="7" heatid="2003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:44.14" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="5259" eventid="6" status="DSQ" swimtime="00:00:51.28" lane="6" heatid="6001" comment="Wechselbeinschläge während der gesamten Schwimmstrecke." />
                <RESULT resultid="5260" eventid="11" swimtime="00:01:32.21" lane="7" heatid="11004" />
                <RESULT resultid="5261" eventid="13" swimtime="00:00:38.79" lane="3" heatid="13003" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1124" birthdate="2011-01-01" gender="M" lastname="Mykhailyk" firstname="Bogdan" license="457896">
              <RESULTS>
                <RESULT resultid="5262" eventid="4" swimtime="00:02:00.14" lane="7" heatid="4003" />
                <RESULT resultid="5263" eventid="6" swimtime="00:00:49.09" lane="2" heatid="6001" />
                <RESULT resultid="5264" eventid="11" swimtime="00:01:42.57" lane="4" heatid="11004" />
                <RESULT resultid="5265" eventid="13" swimtime="00:00:36.07" lane="5" heatid="13009" />
                <RESULT resultid="5266" eventid="24" swimtime="00:03:09.46" lane="1" heatid="24004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:31.87" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="5267" eventid="26" swimtime="00:00:44.95" lane="6" heatid="26017" />
                <RESULT resultid="5268" eventid="34" swimtime="00:01:24.65" lane="3" heatid="34008" />
                <RESULT resultid="5269" eventid="38" swimtime="00:03:42.13" lane="6" heatid="38001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:49.40" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1125" birthdate="2011-01-01" gender="M" lastname="Dreher" firstname="Elias" license="429233">
              <RESULTS>
                <RESULT resultid="5270" eventid="2" swimtime="00:03:15.42" lane="4" heatid="2004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:32.77" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="5271" eventid="4" swimtime="00:01:44.49" lane="4" heatid="4005" />
                <RESULT resultid="5272" eventid="6" swimtime="00:00:40.13" lane="3" heatid="6005" />
                <RESULT resultid="5273" eventid="15" swimtime="00:03:37.81" lane="5" heatid="15003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:45.53" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1126" birthdate="2009-01-01" gender="F" lastname="Thamm" firstname="Elisa" license="397507">
              <RESULTS>
                <RESULT resultid="5274" eventid="23" swimtime="00:02:41.14" lane="5" heatid="23008">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:18.31" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="5275" eventid="25" swimtime="00:00:40.62" lane="2" heatid="25029" />
                <RESULT resultid="5276" eventid="33" swimtime="00:01:10.88" lane="6" heatid="33016" />
                <RESULT resultid="5277" eventid="37" swimtime="00:03:07.75" lane="3" heatid="37005">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:32.65" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1127" birthdate="2011-01-01" gender="F" lastname="Donath" firstname="Emma" license="429234">
              <RESULTS>
                <RESULT resultid="5278" eventid="3" swimtime="00:01:42.18" lane="8" heatid="3008" />
                <RESULT resultid="5279" eventid="5" swimtime="00:00:46.11" lane="4" heatid="5004" />
                <RESULT resultid="5280" eventid="10" swimtime="00:01:35.78" lane="1" heatid="10007" />
                <RESULT resultid="5281" eventid="12" swimtime="00:00:39.44" lane="4" heatid="12004" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1128" birthdate="2011-01-01" gender="M" lastname="Holz" firstname="Florian" license="425562">
              <RESULTS>
                <RESULT resultid="5282" eventid="2" swimtime="00:03:27.40" lane="6" heatid="2004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:40.94" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="5283" eventid="6" swimtime="00:00:43.23" lane="1" heatid="6005" />
                <RESULT resultid="5284" eventid="11" swimtime="00:01:36.67" lane="2" heatid="11007" />
                <RESULT resultid="5285" eventid="13" swimtime="00:00:36.47" lane="5" heatid="13008" />
                <RESULT resultid="5286" eventid="24" status="DNS" swimtime="00:00:00.00" lane="3" heatid="24005" />
                <RESULT resultid="5287" eventid="26" status="DNS" swimtime="00:00:00.00" lane="3" heatid="26018" />
                <RESULT resultid="5288" eventid="34" status="DNS" swimtime="00:00:00.00" lane="3" heatid="34009" />
                <RESULT resultid="5289" eventid="38" status="DNS" swimtime="00:00:00.00" lane="1" heatid="38003" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1129" birthdate="2014-01-01" gender="F" lastname="Thomas" firstname="Fritzi" license="451398">
              <RESULTS>
                <RESULT resultid="5290" eventid="19" swimtime="00:00:56.52" lane="6" heatid="19003" />
                <RESULT resultid="5291" eventid="21" swimtime="00:01:10.03" lane="8" heatid="21004" />
                <RESULT resultid="5292" eventid="25" swimtime="00:00:53.71" lane="1" heatid="25006" />
                <RESULT resultid="5293" eventid="29" swimtime="00:00:45.37" lane="7" heatid="29003" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1130" birthdate="2008-01-01" gender="F" lastname="Prill" firstname="Isabell" license="378819">
              <RESULTS>
                <RESULT resultid="5294" eventid="19" swimtime="00:00:49.45" lane="1" heatid="19022" />
                <RESULT resultid="5295" eventid="25" swimtime="00:00:40.61" lane="5" heatid="25029" />
                <RESULT resultid="5296" eventid="33" swimtime="00:01:24.01" lane="2" heatid="33010" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1131" birthdate="2011-01-01" gender="F" lastname="Gunsilius" firstname="Jette" license="425560">
              <RESULTS>
                <RESULT resultid="5297" eventid="23" swimtime="00:02:41.25" lane="2" heatid="23008">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:17.16" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="5298" eventid="25" swimtime="00:00:39.21" lane="8" heatid="25030" />
                <RESULT resultid="5299" eventid="33" swimtime="00:01:12.66" lane="5" heatid="33013" />
                <RESULT resultid="5300" eventid="37" swimtime="00:03:01.38" lane="6" heatid="37005">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:27.74" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1132" birthdate="2012-01-01" gender="F" lastname="Menzel" firstname="Jette" license="442930">
              <RESULTS>
                <RESULT resultid="5301" eventid="19" status="DNS" swimtime="00:00:00.00" lane="5" heatid="19012" />
                <RESULT resultid="5302" eventid="23" status="DNS" swimtime="00:00:00.00" lane="6" heatid="23004" />
                <RESULT resultid="5303" eventid="25" status="DNS" swimtime="00:00:00.00" lane="2" heatid="25007" />
                <RESULT resultid="5304" eventid="33" status="DNS" swimtime="00:00:00.00" lane="3" heatid="33007" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1133" birthdate="2012-01-01" gender="M" lastname="Bormann" firstname="Julian" license="442932">
              <RESULTS>
                <RESULT resultid="5305" eventid="4" swimtime="00:01:40.44" lane="6" heatid="4006" />
                <RESULT resultid="5306" eventid="11" swimtime="00:01:38.54" lane="4" heatid="11002" />
                <RESULT resultid="5307" eventid="13" swimtime="00:00:37.21" lane="7" heatid="13003" />
                <RESULT resultid="5308" eventid="15" swimtime="00:03:43.75" lane="5" heatid="15004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:48.77" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="5309" eventid="20" swimtime="00:00:46.65" lane="8" heatid="20016" />
                <RESULT resultid="5310" eventid="26" swimtime="00:00:46.82" lane="7" heatid="26014" />
                <RESULT resultid="5311" eventid="36" swimtime="00:01:51.73" lane="3" heatid="36001" />
                <RESULT resultid="5312" eventid="38" swimtime="00:03:30.70" lane="2" heatid="38001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:44.27" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1134" birthdate="2007-01-01" gender="M" lastname="Simon" firstname="Julius" license="356385">
              <RESULTS>
                <RESULT resultid="5313" eventid="2" swimtime="00:02:34.46" lane="7" heatid="2008">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:08.86" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="5314" eventid="11" swimtime="00:01:06.85" lane="4" heatid="11012" />
                <RESULT resultid="5315" eventid="13" swimtime="00:00:26.17" lane="1" heatid="13018" />
                <RESULT resultid="5316" eventid="26" swimtime="00:00:29.77" lane="5" heatid="26024" />
                <RESULT resultid="5317" eventid="34" swimtime="00:00:58.44" lane="4" heatid="34014" />
                <RESULT resultid="5318" eventid="38" swimtime="00:02:28.35" lane="3" heatid="38005">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:11.95" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1135" birthdate="2009-01-01" gender="F" lastname="Fornfeist" firstname="Kiara" license="397503">
              <RESULTS>
                <RESULT resultid="5319" eventid="3" swimtime="00:01:43.54" lane="1" heatid="3008" />
                <RESULT resultid="5320" eventid="5" swimtime="00:00:37.92" lane="6" heatid="5010" />
                <RESULT resultid="5321" eventid="10" swimtime="00:01:27.44" lane="1" heatid="10013" />
                <RESULT resultid="5322" eventid="19" status="DNS" swimtime="00:00:00.00" lane="7" heatid="19023" />
                <RESULT resultid="5323" eventid="25" status="DNS" swimtime="00:00:00.00" lane="4" heatid="25030" />
                <RESULT resultid="5324" eventid="35" status="DNS" swimtime="00:00:00.00" lane="1" heatid="35003" />
                <RESULT resultid="5325" eventid="37" status="DNS" swimtime="00:00:00.00" lane="4" heatid="37006" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1136" birthdate="2010-01-01" gender="F" lastname="Saremsky" firstname="Lisa" license="415165">
              <RESULTS>
                <RESULT resultid="5326" eventid="1" swimtime="00:03:10.81" lane="5" heatid="1004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:29.14" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="5327" eventid="5" swimtime="00:00:36.85" lane="1" heatid="5011" />
                <RESULT resultid="5328" eventid="10" swimtime="00:01:27.16" lane="5" heatid="10012" />
                <RESULT resultid="5329" eventid="25" status="DNS" swimtime="00:00:00.00" lane="8" heatid="25031" />
                <RESULT resultid="5330" eventid="37" status="DNS" swimtime="00:00:00.00" lane="5" heatid="37005" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1137" birthdate="2009-01-01" gender="F" lastname="Gunsilius" firstname="Luisa" license="397501">
              <RESULTS>
                <RESULT resultid="5331" eventid="23" swimtime="00:02:41.59" lane="4" heatid="23008">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:17.34" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="5332" eventid="25" swimtime="00:00:38.24" lane="5" heatid="25031" />
                <RESULT resultid="5333" eventid="33" swimtime="00:01:11.82" lane="3" heatid="33015" />
                <RESULT resultid="5334" eventid="37" swimtime="00:02:55.35" lane="5" heatid="37006">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:25.22" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1138" birthdate="2013-01-01" gender="M" lastname="Nowotny" firstname="Lukas" license="445777">
              <RESULTS>
                <RESULT resultid="5335" eventid="2" swimtime="00:03:43.43" lane="6" heatid="2002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:45.71" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="5336" eventid="6" swimtime="00:00:50.77" lane="4" heatid="6001" />
                <RESULT resultid="5337" eventid="13" swimtime="00:00:41.64" lane="5" heatid="13001" />
                <RESULT resultid="5338" eventid="15" swimtime="00:04:12.83" lane="5" heatid="15002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:02:02.03" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1139" birthdate="2012-01-01" gender="F" lastname="Illing" firstname="Lynn Xenia" license="436674">
              <RESULTS>
                <RESULT resultid="5339" eventid="1" swimtime="00:02:55.98" lane="1" heatid="1007">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:24.53" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="5340" eventid="3" swimtime="00:01:31.09" lane="3" heatid="3010" />
                <RESULT resultid="5341" eventid="5" swimtime="00:00:35.34" lane="8" heatid="5012" />
                <RESULT resultid="5342" eventid="10" swimtime="00:01:21.13" lane="8" heatid="10015" />
                <RESULT resultid="5343" eventid="17" swimtime="00:00:44.70" lane="4" heatid="17016" />
                <RESULT resultid="5344" eventid="25" swimtime="00:00:36.82" lane="8" heatid="25033" />
                <RESULT resultid="5345" eventid="31" swimtime="00:00:42.95" lane="4" heatid="31007" />
                <RESULT resultid="5346" eventid="35" swimtime="00:01:22.72" lane="8" heatid="35004" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1140" birthdate="2012-01-01" gender="F" lastname="Tschirner" firstname="Marah" license="442928">
              <RESULTS>
                <RESULT resultid="5347" eventid="1" status="WDR" swimtime="00:00:00.00" lane="8" heatid="1003" />
                <RESULT resultid="5348" eventid="5" status="WDR" swimtime="00:00:00.00" lane="2" heatid="5006" />
                <RESULT resultid="5349" eventid="10" status="WDR" swimtime="00:00:00.00" lane="1" heatid="10004" />
                <RESULT resultid="5350" eventid="12" status="WDR" swimtime="00:00:00.00" lane="4" heatid="12009" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1141" birthdate="2009-01-01" gender="F" lastname="Thamm" firstname="Marie" license="397505">
              <RESULTS>
                <RESULT resultid="5351" eventid="1" swimtime="00:02:50.45" lane="6" heatid="1006">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:20.37" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="5352" eventid="5" swimtime="00:00:32.97" lane="6" heatid="5013" />
                <RESULT resultid="5353" eventid="10" swimtime="00:01:18.82" lane="2" heatid="10015" />
                <RESULT resultid="5354" eventid="12" swimtime="00:00:29.72" lane="7" heatid="12018" />
                <RESULT resultid="5355" eventid="23" swimtime="00:02:30.47" lane="2" heatid="23010">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:12.17" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="5356" eventid="25" swimtime="00:00:35.62" lane="8" heatid="25034" />
                <RESULT resultid="5357" eventid="33" swimtime="00:01:05.45" lane="3" heatid="33018" />
                <RESULT resultid="5358" eventid="35" swimtime="00:01:16.20" lane="5" heatid="35004" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1142" birthdate="2008-01-01" gender="M" lastname="Woite" firstname="Miko" license="354185">
              <RESULTS>
                <RESULT resultid="5359" eventid="4" swimtime="00:01:23.85" lane="4" heatid="4010" />
                <RESULT resultid="5360" eventid="6" swimtime="00:00:30.85" lane="4" heatid="6010" />
                <RESULT resultid="5361" eventid="15" swimtime="00:03:03.35" lane="8" heatid="15007">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:26.65" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="5362" eventid="20" swimtime="00:00:37.28" lane="3" heatid="20021" />
                <RESULT resultid="5363" eventid="24" swimtime="00:02:21.71" lane="2" heatid="24009">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:08.17" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="5364" eventid="36" swimtime="00:01:11.33" lane="6" heatid="36003" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1143" birthdate="2010-01-01" gender="F" lastname="Woite" firstname="Mira" license="415160">
              <RESULTS>
                <RESULT resultid="5365" eventid="1" swimtime="00:03:29.39" lane="6" heatid="1002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:37.51" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="5366" eventid="3" swimtime="00:01:46.48" lane="5" heatid="3007" />
                <RESULT resultid="5367" eventid="5" swimtime="00:00:41.31" lane="1" heatid="5008" />
                <RESULT resultid="5369" eventid="14" swimtime="00:03:36.05" lane="4" heatid="14004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:47.02" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="5370" eventid="19" swimtime="00:00:48.82" lane="1" heatid="19020" />
                <RESULT resultid="5371" eventid="25" swimtime="00:00:45.42" lane="4" heatid="25019" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1144" birthdate="2007-01-01" gender="M" lastname="Saremsky" firstname="Moritz" license="363799">
              <RESULTS>
                <RESULT resultid="5372" eventid="20" swimtime="00:00:36.68" lane="6" heatid="20022" />
                <RESULT resultid="5373" eventid="26" swimtime="00:00:36.09" lane="4" heatid="26022" />
                <RESULT resultid="5374" eventid="34" swimtime="00:01:07.94" lane="8" heatid="34013" />
                <RESULT resultid="5375" eventid="36" swimtime="00:01:16.88" lane="1" heatid="36003" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1145" birthdate="2014-01-01" gender="F" lastname="Petersohn" firstname="Nele Kristin" license="451396">
              <RESULTS>
                <RESULT resultid="5376" eventid="19" swimtime="00:00:50.35" lane="5" heatid="19018" />
                <RESULT resultid="5377" eventid="25" swimtime="00:00:46.87" lane="5" heatid="25019" />
                <RESULT resultid="5378" eventid="27" swimtime="00:01:02.28" lane="6" heatid="27005" />
                <RESULT resultid="5379" eventid="29" swimtime="00:00:42.37" lane="5" heatid="29012" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1146" birthdate="2014-01-01" gender="F" lastname="Eifler" firstname="Nelly" license="451392">
              <RESULTS>
                <RESULT resultid="5380" eventid="19" swimtime="00:00:53.26" lane="7" heatid="19013" />
                <RESULT resultid="5381" eventid="21" swimtime="00:00:57.15" lane="7" heatid="21011" />
                <RESULT resultid="5382" eventid="25" status="DSQ" swimtime="00:00:46.09" lane="7" heatid="25022" comment="Der Zielanschlag erfolgte nich in Rückenlage." />
                <RESULT resultid="5383" eventid="29" swimtime="00:00:40.01" lane="7" heatid="29013" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1147" birthdate="2008-01-01" gender="M" lastname="Nitsche" firstname="Niklas" license="378824">
              <RESULTS>
                <RESULT resultid="5384" eventid="2" swimtime="00:02:49.86" lane="3" heatid="2006">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:18.64" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="5385" eventid="6" swimtime="00:00:33.66" lane="3" heatid="6008" />
                <RESULT resultid="5386" eventid="11" swimtime="00:01:16.55" lane="6" heatid="11011" />
                <RESULT resultid="5387" eventid="26" swimtime="00:00:34.06" lane="6" heatid="26023" />
                <RESULT resultid="5388" eventid="38" swimtime="00:02:46.41" lane="4" heatid="38004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:18.78" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1148" birthdate="2010-01-01" gender="F" lastname="Pleschinger" firstname="Penelope" license="399989">
              <RESULTS>
                <RESULT resultid="5389" eventid="3" swimtime="00:01:29.74" lane="4" heatid="3010" />
                <RESULT resultid="5390" eventid="5" swimtime="00:00:35.25" lane="3" heatid="5013" />
                <RESULT resultid="5391" eventid="10" swimtime="00:01:16.53" lane="2" heatid="10016" />
                <RESULT resultid="5392" eventid="14" swimtime="00:03:11.77" lane="1" heatid="14007">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:33.27" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="5393" eventid="23" swimtime="00:02:30.32" lane="2" heatid="23011">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:10.48" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="5394" eventid="25" swimtime="00:00:34.88" lane="1" heatid="25034" />
                <RESULT resultid="5395" eventid="37" swimtime="00:02:46.46" lane="5" heatid="37007">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:21.88" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1149" birthdate="2014-01-01" gender="F" lastname="Dreher" firstname="Rosalie" license="451391">
              <RESULTS>
                <RESULT resultid="5396" eventid="17" swimtime="00:01:08.45" lane="8" heatid="17004" />
                <RESULT resultid="5397" eventid="19" swimtime="00:00:56.57" lane="4" heatid="19008" />
                <RESULT resultid="5398" eventid="25" swimtime="00:00:52.09" lane="2" heatid="25014" />
                <RESULT resultid="5399" eventid="29" swimtime="00:00:48.65" lane="7" heatid="29007" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1150" birthdate="2011-01-01" gender="F" lastname="Petersohn" firstname="Sophie Marie" license="434411">
              <RESULTS>
                <RESULT resultid="5400" eventid="1" swimtime="00:03:02.44" lane="2" heatid="1004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:27.71" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="5401" eventid="3" swimtime="00:01:34.77" lane="1" heatid="3009" />
                <RESULT resultid="5402" eventid="5" swimtime="00:00:36.90" lane="3" heatid="5010" />
                <RESULT resultid="5403" eventid="10" swimtime="00:01:30.07" lane="1" heatid="10012" />
                <RESULT resultid="5404" eventid="19" swimtime="00:00:43.01" lane="4" heatid="19024" />
                <RESULT resultid="5405" eventid="25" swimtime="00:00:37.60" lane="4" heatid="25023" />
                <RESULT resultid="5406" eventid="35" swimtime="00:01:20.74" lane="4" heatid="35003" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1151" birthdate="2014-01-01" gender="M" lastname="Steinert" firstname="Tom Raphael" license="451401">
              <RESULTS>
                <RESULT resultid="5407" eventid="20" swimtime="00:00:53.67" lane="3" heatid="20007" />
                <RESULT resultid="5408" eventid="26" swimtime="00:00:50.34" lane="1" heatid="26008" />
                <RESULT resultid="5409" eventid="28" swimtime="00:01:04.00" lane="7" heatid="28006" />
                <RESULT resultid="5410" eventid="30" swimtime="00:00:51.17" lane="5" heatid="30004" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1152" birthdate="2012-01-01" gender="M" lastname="Steudtner" firstname="Vincent" license="442934">
              <RESULTS>
                <RESULT resultid="5411" eventid="2" status="DNS" swimtime="00:00:00.00" lane="6" heatid="2005" />
                <RESULT resultid="5412" eventid="6" swimtime="00:00:41.46" lane="8" heatid="6007" />
                <RESULT resultid="5413" eventid="11" status="DNS" swimtime="00:00:00.00" lane="3" heatid="11008" />
                <RESULT resultid="5414" eventid="13" swimtime="00:00:32.44" lane="5" heatid="13012" />
                <RESULT resultid="5415" eventid="20" status="DNS" swimtime="00:00:00.00" lane="4" heatid="20018" />
                <RESULT resultid="5416" eventid="26" status="DNS" swimtime="00:00:00.00" lane="1" heatid="26020" />
                <RESULT resultid="5417" eventid="34" status="DNS" swimtime="00:00:00.00" lane="3" heatid="34012" />
                <RESULT resultid="5418" eventid="38" status="DNS" swimtime="00:00:00.00" lane="3" heatid="38003" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY number="1" gender="X" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="5251" eventid="16" swimtime="00:02:09.89" lane="3" heatid="16002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:08.13" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1134" number="1" />
                    <RELAYPOSITION athleteid="1142" number="2" />
                    <RELAYPOSITION athleteid="1141" number="3" />
                    <RELAYPOSITION athleteid="1147" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" gender="X" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="5252" eventid="7" swimtime="00:02:25.72" lane="2" heatid="7003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:18.75" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1148" number="1" />
                    <RELAYPOSITION athleteid="1152" number="2" />
                    <RELAYPOSITION athleteid="1139" number="3" />
                    <RELAYPOSITION athleteid="1122" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="2" gender="X" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="5253" eventid="7" swimtime="00:02:30.88" lane="4" heatid="7002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:22.11" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1136" number="1" />
                    <RELAYPOSITION athleteid="1133" number="2" />
                    <RELAYPOSITION athleteid="1150" number="3" />
                    <RELAYPOSITION athleteid="1125" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="3" gender="X" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="5254" eventid="7" swimtime="00:02:43.72" lane="6" heatid="7002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:27.63" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1128" number="1" />
                    <RELAYPOSITION athleteid="1127" number="2" />
                    <RELAYPOSITION athleteid="1143" number="3" />
                    <RELAYPOSITION athleteid="1124" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB name="SV Lok Leipzig-Mitte e.V." nation="GER" region="12" code="3393">
          <ATHLETES>
            <ATHLETE athleteid="720" birthdate="2013-01-01" gender="M" lastname="Brauer" firstname="Fabian" license="445392">
              <RESULTS>
                <RESULT resultid="3439" eventid="6" swimtime="00:00:38.12" lane="5" heatid="6006" />
                <RESULT resultid="3438" eventid="11" swimtime="00:01:32.15" lane="7" heatid="11008" />
                <RESULT resultid="3437" eventid="13" swimtime="00:00:33.04" lane="2" heatid="13012" />
                <RESULT resultid="3436" eventid="22" swimtime="00:00:44.40" lane="5" heatid="22011" />
                <RESULT resultid="3435" eventid="24" swimtime="00:02:45.58" lane="1" heatid="24006">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:22.60" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="3434" eventid="34" swimtime="00:01:14.94" lane="2" heatid="34011" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="SV Weixdorf e.V." nation="GER" region="12" code="3366">
          <ATHLETES>
            <ATHLETE athleteid="35" birthdate="2015-01-01" gender="M" lastname="Jahn" firstname="Anton" license="448908">
              <RESULTS>
                <RESULT resultid="193" eventid="18" swimtime="00:01:17.68" lane="8" heatid="18004" />
                <RESULT resultid="194" eventid="22" swimtime="00:01:13.48" lane="7" heatid="22002" />
                <RESULT resultid="195" eventid="26" swimtime="00:01:05.88" lane="4" heatid="26001" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="36" birthdate="2015-01-01" gender="F" lastname="Witt" firstname="Aria Luise" license="467915">
              <RESULTS>
                <RESULT resultid="197" eventid="17" swimtime="00:01:02.68" lane="1" heatid="17005" />
                <RESULT resultid="198" eventid="21" swimtime="00:01:03.73" lane="8" heatid="21007" />
                <RESULT resultid="199" eventid="25" swimtime="00:00:52.52" lane="1" heatid="25010" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="37" birthdate="2012-01-01" gender="M" lastname="Marschner" firstname="Ben" license="448906">
              <RESULTS>
                <RESULT resultid="201" eventid="18" swimtime="00:00:58.45" lane="1" heatid="18010" />
                <RESULT resultid="202" eventid="20" swimtime="00:01:09.75" lane="2" heatid="20002" />
                <RESULT resultid="203" eventid="26" swimtime="00:00:51.43" lane="3" heatid="26009" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="38" birthdate="2015-01-01" gender="M" lastname="Juen" firstname="Darian" license="448909">
              <RESULTS>
                <RESULT resultid="204" eventid="18" swimtime="00:01:10.95" lane="6" heatid="18003" />
                <RESULT resultid="205" eventid="22" swimtime="00:01:07.75" lane="2" heatid="22003" />
                <RESULT resultid="206" eventid="26" swimtime="00:00:59.33" lane="4" heatid="26004" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="39" birthdate="2013-01-01" gender="F" lastname="Koenig" firstname="Dorothea" license="424080">
              <RESULTS>
                <RESULT resultid="208" eventid="10" swimtime="00:01:34.79" lane="3" heatid="10007" />
                <RESULT resultid="209" eventid="12" swimtime="00:00:35.69" lane="2" heatid="12009" />
                <RESULT resultid="210" eventid="14" swimtime="00:03:51.76" lane="8" heatid="14003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:52.13" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="211" eventid="19" swimtime="00:00:48.13" lane="6" heatid="19016" />
                <RESULT resultid="212" eventid="23" swimtime="00:03:08.79" lane="4" heatid="23003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:28.85" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="213" eventid="25" swimtime="00:00:42.67" lane="5" heatid="25024" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="40" birthdate="2015-01-01" gender="M" lastname="Hickmann" firstname="Finjas" license="459062">
              <RESULTS>
                <RESULT resultid="215" eventid="18" swimtime="00:01:13.97" lane="7" heatid="18003" />
                <RESULT resultid="216" eventid="22" swimtime="00:01:15.56" lane="5" heatid="22001" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="41" birthdate="2011-01-01" gender="F" lastname="Buder" firstname="Freya" license="397759">
              <RESULTS>
                <RESULT resultid="218" eventid="10" swimtime="00:01:24.70" lane="8" heatid="10012" />
                <RESULT resultid="219" eventid="37" swimtime="00:02:57.51" lane="3" heatid="37006">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:27.64" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="42" birthdate="2015-01-01" gender="F" lastname="Czarnecki" firstname="Greta Luise" license="448905">
              <RESULTS>
                <RESULT resultid="220" eventid="19" swimtime="00:01:00.66" lane="3" heatid="19004" />
                <RESULT resultid="221" eventid="21" swimtime="00:01:15.65" lane="2" heatid="21005" />
                <RESULT resultid="222" eventid="25" swimtime="00:00:52.91" lane="1" heatid="25015" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="43" birthdate="2011-01-01" gender="F" lastname="Riedel" firstname="Hilda" license="412725">
              <RESULTS>
                <RESULT resultid="224" eventid="19" swimtime="00:00:53.76" lane="2" heatid="19013" />
                <RESULT resultid="225" eventid="23" swimtime="00:03:13.55" lane="8" heatid="23003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:35.72" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="226" eventid="25" swimtime="00:00:45.06" lane="2" heatid="25021" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="44" birthdate="2014-01-01" gender="F" lastname="Schuster" firstname="Leonie" license="448904">
              <RESULTS>
                <RESULT resultid="227" eventid="17" swimtime="00:01:09.07" lane="2" heatid="17006" />
                <RESULT resultid="228" eventid="21" swimtime="00:01:15.21" lane="4" heatid="21003" />
                <RESULT resultid="229" eventid="25" swimtime="00:01:00.71" lane="3" heatid="25009" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="45" birthdate="2009-01-01" gender="M" lastname="Pfützner" firstname="Matteo" license="397752">
              <RESULTS>
                <RESULT resultid="231" eventid="11" swimtime="00:01:35.71" lane="3" heatid="11003" />
                <RESULT resultid="232" eventid="13" status="DSQ" swimtime="00:00:31.36" lane="1" heatid="13013" comment="Start vor dem Startsignal." />
                <RESULT resultid="233" eventid="15" swimtime="00:03:37.39" lane="8" heatid="15006">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:38.85" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="46" birthdate="2010-01-01" gender="F" lastname="Albrecht" firstname="Mia" license="404147">
              <RESULTS>
                <RESULT resultid="234" eventid="3" swimtime="00:01:21.82" lane="4" heatid="3011" />
                <RESULT resultid="235" eventid="8" swimtime="00:02:35.92" lane="4" heatid="8001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:13.53" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="47" birthdate="2014-01-01" gender="M" lastname="Marschner" firstname="Oskar" license="448907">
              <RESULTS>
                <RESULT resultid="236" eventid="18" swimtime="00:01:14.09" lane="2" heatid="18006" />
                <RESULT resultid="237" eventid="22" swimtime="00:01:09.71" lane="5" heatid="22002" />
                <RESULT resultid="238" eventid="26" swimtime="00:00:53.94" lane="6" heatid="26007" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="48" birthdate="2010-01-01" gender="M" lastname="Liepke" firstname="Paul" license="397757">
              <RESULTS>
                <RESULT resultid="240" eventid="4" swimtime="00:01:15.23" lane="5" heatid="4011" />
                <RESULT resultid="241" eventid="9" swimtime="00:02:39.75" lane="3" heatid="9001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:17.40" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="49" birthdate="2013-01-01" gender="F" lastname="Liepke" firstname="Thea" license="424069">
              <RESULTS>
                <RESULT resultid="242" eventid="10" swimtime="00:01:33.57" lane="8" heatid="10008" />
                <RESULT resultid="243" eventid="12" swimtime="00:00:38.14" lane="8" heatid="12005" />
                <RESULT resultid="244" eventid="14" swimtime="00:03:58.66" lane="3" heatid="14002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:56.70" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="245" eventid="19" swimtime="00:00:53.33" lane="1" heatid="19011" />
                <RESULT resultid="246" eventid="23" swimtime="00:03:07.58" lane="7" heatid="23003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:31.97" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="247" eventid="25" swimtime="00:00:43.83" lane="8" heatid="25023" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="SV Zwickau von 1904" nation="GER" region="12" code="3400">
          <ATHLETES>
            <ATHLETE athleteid="1106" birthdate="2014-01-01" gender="M" lastname="Plettig" firstname="Ben" license="464151">
              <RESULTS>
                <RESULT resultid="5183" eventid="18" swimtime="00:01:10.36" lane="6" heatid="18005" />
                <RESULT resultid="5184" eventid="20" swimtime="00:01:03.12" lane="8" heatid="20004" />
                <RESULT resultid="5185" eventid="26" swimtime="00:00:50.02" lane="8" heatid="26009" />
                <RESULT resultid="5186" eventid="30" swimtime="00:00:47.92" lane="3" heatid="30004" />
                <RESULT resultid="5187" eventid="34" swimtime="00:01:51.32" lane="3" heatid="34001" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1107" birthdate="2013-01-01" gender="F" lastname="Dressel" firstname="Clara" license="447504">
              <RESULTS>
                <RESULT resultid="5188" eventid="1" swimtime="00:03:48.46" lane="5" heatid="1001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:50.12" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="5189" eventid="5" swimtime="00:00:55.63" lane="3" heatid="5001" />
                <RESULT resultid="5190" eventid="10" swimtime="00:01:42.39" lane="8" heatid="10004" />
                <RESULT resultid="5191" eventid="12" swimtime="00:00:41.00" lane="6" heatid="12003" />
                <RESULT resultid="5192" eventid="23" swimtime="00:03:16.26" lane="3" heatid="23002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:34.97" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="5193" eventid="25" swimtime="00:00:48.01" lane="6" heatid="25017" />
                <RESULT resultid="5194" eventid="33" swimtime="00:01:30.32" lane="3" heatid="33005" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1108" birthdate="2014-01-01" gender="M" lastname="Zänsler" firstname="Elias" license="461989">
              <RESULTS>
                <RESULT resultid="5195" eventid="18" swimtime="00:01:16.47" lane="2" heatid="18004" />
                <RESULT resultid="5196" eventid="20" swimtime="00:01:03.98" lane="3" heatid="20002" />
                <RESULT resultid="5197" eventid="26" swimtime="00:00:54.70" lane="2" heatid="26004" />
                <RESULT resultid="5198" eventid="30" swimtime="00:00:53.45" lane="7" heatid="30002" />
                <RESULT resultid="5199" eventid="32" swimtime="00:01:09.51" lane="3" heatid="32002" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1109" birthdate="2015-01-01" gender="F" lastname="Birzer" firstname="Frieda" license="466284">
              <RESULTS>
                <RESULT resultid="5200" eventid="17" swimtime="00:01:12.06" lane="4" heatid="17006" />
                <RESULT resultid="5201" eventid="19" swimtime="00:00:56.98" lane="5" heatid="19009" />
                <RESULT resultid="5202" eventid="25" swimtime="00:00:54.52" lane="2" heatid="25008" />
                <RESULT resultid="5203" eventid="27" swimtime="00:01:04.57" lane="7" heatid="27001" />
                <RESULT resultid="5204" eventid="29" swimtime="00:00:51.17" lane="4" heatid="29006" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1110" birthdate="2010-01-01" gender="F" lastname="Flemming" firstname="Heda" license="410490">
              <RESULTS>
                <RESULT resultid="5205" eventid="3" swimtime="00:01:36.73" lane="6" heatid="3010" />
                <RESULT resultid="5206" eventid="5" swimtime="00:00:37.77" lane="8" heatid="5010" />
                <RESULT resultid="5207" eventid="10" swimtime="00:01:22.42" lane="8" heatid="10014" />
                <RESULT resultid="5208" eventid="12" swimtime="00:00:34.25" lane="6" heatid="12016" />
                <RESULT resultid="5209" eventid="19" swimtime="00:00:42.92" lane="4" heatid="19025" />
                <RESULT resultid="5210" eventid="25" swimtime="00:00:37.87" lane="4" heatid="25033" />
                <RESULT resultid="5211" eventid="33" swimtime="00:01:16.71" lane="4" heatid="33014" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1111" birthdate="2014-01-01" gender="F" lastname="Sprenger" firstname="Lara" license="456271">
              <RESULTS>
                <RESULT resultid="5212" eventid="17" swimtime="00:00:57.56" lane="7" heatid="17014" />
                <RESULT resultid="5213" eventid="21" swimtime="00:01:00.74" lane="2" heatid="21010" />
                <RESULT resultid="5214" eventid="25" swimtime="00:00:48.13" lane="7" heatid="25018" />
                <RESULT resultid="5215" eventid="29" swimtime="00:00:42.33" lane="5" heatid="29010" />
                <RESULT resultid="5216" eventid="31" swimtime="00:01:10.27" lane="8" heatid="31003" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1112" birthdate="2013-01-01" gender="F" lastname="Schneider" firstname="Laura" license="447503">
              <RESULTS>
                <RESULT resultid="5217" eventid="3" swimtime="00:01:37.49" lane="6" heatid="3006" />
                <RESULT resultid="5218" eventid="5" swimtime="00:00:42.89" lane="1" heatid="5006" />
                <RESULT resultid="5219" eventid="10" swimtime="00:01:34.07" lane="8" heatid="10009" />
                <RESULT resultid="5220" eventid="14" swimtime="00:03:45.44" lane="8" heatid="14004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:47.46" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="5221" eventid="19" swimtime="00:00:44.37" lane="7" heatid="19021" />
                <RESULT resultid="5222" eventid="21" swimtime="00:00:52.20" lane="2" heatid="21012" />
                <RESULT resultid="5223" eventid="25" swimtime="00:00:42.00" lane="6" heatid="25029" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1113" birthdate="2015-01-01" gender="F" lastname="Schneider" firstname="Linda" license="466281">
              <RESULTS>
                <RESULT resultid="5224" eventid="19" swimtime="00:01:01.61" lane="3" heatid="19002" />
                <RESULT resultid="5225" eventid="21" swimtime="00:01:06.26" lane="4" heatid="21005" />
                <RESULT resultid="5226" eventid="25" swimtime="00:00:56.22" lane="2" heatid="25003" />
                <RESULT resultid="5227" eventid="29" swimtime="00:00:55.02" lane="2" heatid="29002" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1114" birthdate="2012-01-01" gender="F" lastname="Komar" firstname="Lindsay" license="436924">
              <RESULTS>
                <RESULT resultid="5228" eventid="1" swimtime="00:03:18.27" lane="7" heatid="1004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:34.97" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="5229" eventid="5" swimtime="00:00:38.77" lane="1" heatid="5009" />
                <RESULT resultid="5230" eventid="8" swimtime="00:03:34.45" lane="2" heatid="8001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:37.20" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="5231" eventid="12" swimtime="00:00:35.78" lane="1" heatid="12012" />
                <RESULT resultid="5232" eventid="19" swimtime="00:00:46.53" lane="2" heatid="19021" />
                <RESULT resultid="5233" eventid="25" swimtime="00:00:40.70" lane="2" heatid="25026" />
                <RESULT resultid="5234" eventid="31" swimtime="00:00:59.39" lane="6" heatid="31005" />
                <RESULT resultid="5235" eventid="35" swimtime="00:01:34.13" lane="5" heatid="35002" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1115" birthdate="2010-01-01" gender="F" lastname="Rohatzsch" firstname="Maxime" license="410491">
              <RESULTS>
                <RESULT resultid="5236" eventid="1" swimtime="00:02:59.68" lane="2" heatid="1005">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:23.79" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="5237" eventid="5" swimtime="00:00:36.80" lane="2" heatid="5008" />
                <RESULT resultid="5238" eventid="10" swimtime="00:01:20.67" lane="4" heatid="10014" />
                <RESULT resultid="5239" eventid="12" swimtime="00:00:32.44" lane="2" heatid="12015" />
                <RESULT resultid="5240" eventid="23" swimtime="00:02:35.93" lane="5" heatid="23010">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:15.07" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="5241" eventid="25" swimtime="00:00:37.33" lane="7" heatid="25033" />
                <RESULT resultid="5242" eventid="33" swimtime="00:01:11.39" lane="5" heatid="33016" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1116" birthdate="2010-01-01" gender="M" lastname="Käser" firstname="Mika Marco" license="423052">
              <RESULTS>
                <RESULT resultid="5243" eventid="20" swimtime="00:00:43.31" lane="3" heatid="20018" />
                <RESULT resultid="5244" eventid="24" swimtime="00:02:42.23" lane="7" heatid="24006">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:20.59" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="5245" eventid="26" swimtime="00:00:39.53" lane="2" heatid="26019" />
                <RESULT resultid="5246" eventid="34" swimtime="00:01:13.23" lane="4" heatid="34010" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1117" birthdate="2013-01-01" gender="F" lastname="Zaiaieva" firstname="Vlada" license="468008">
              <RESULTS>
                <RESULT resultid="5247" eventid="17" status="DSQ" swimtime="00:01:06.75" lane="7" heatid="17009" comment="Die Hände wurden während der Schwimmstrecke nicht übereinander gelegt." />
                <RESULT resultid="5248" eventid="21" status="DSQ" swimtime="00:01:04.42" lane="5" heatid="21005" comment="Das Brett wurde beim Anschlag vorn nicht umfasst." />
                <RESULT resultid="5249" eventid="25" swimtime="00:00:50.16" lane="4" heatid="25012" />
                <RESULT resultid="5250" eventid="33" swimtime="00:01:37.76" lane="1" heatid="33004" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="SVV Plauen" nation="GER" region="12" code="6253">
          <ATHLETES>
            <ATHLETE athleteid="1009" birthdate="2015-01-01" gender="M" lastname="Drbal" firstname="Dean" license="471975">
              <RESULTS>
                <RESULT resultid="4679" eventid="18" swimtime="00:01:07.15" lane="7" heatid="18007" />
                <RESULT resultid="4680" eventid="22" swimtime="00:01:09.80" lane="2" heatid="22006" />
                <RESULT resultid="4681" eventid="26" swimtime="00:00:56.08" lane="7" heatid="26006" />
                <RESULT resultid="4682" eventid="30" swimtime="00:00:55.54" lane="1" heatid="30002" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1010" birthdate="2012-01-01" gender="M" lastname="Mocker" firstname="Felix" license="439927">
              <RESULTS>
                <RESULT resultid="4683" eventid="4" status="DNS" swimtime="00:00:00.00" lane="4" heatid="4008" />
                <RESULT resultid="4684" eventid="6" status="DNS" swimtime="00:00:00.00" lane="3" heatid="6006" />
                <RESULT resultid="4685" eventid="15" status="DNS" swimtime="00:00:00.00" lane="6" heatid="15005" />
                <RESULT resultid="4686" eventid="20" status="DNS" swimtime="00:00:00.00" lane="7" heatid="20015" />
                <RESULT resultid="4687" eventid="24" status="DNS" swimtime="00:00:00.00" lane="3" heatid="24006" />
                <RESULT resultid="4688" eventid="28" status="DNS" swimtime="00:00:00.00" lane="3" heatid="28008" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1011" birthdate="2013-01-01" gender="F" lastname="Wunderlich" firstname="Frida-Malin" license="449330">
              <RESULTS>
                <RESULT resultid="4689" eventid="5" swimtime="00:00:55.00" lane="7" heatid="5002" />
                <RESULT resultid="4690" eventid="12" swimtime="00:00:41.17" lane="3" heatid="12004" />
                <RESULT resultid="4691" eventid="14" swimtime="00:04:22.14" lane="7" heatid="14002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:02:07.78" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="4692" eventid="21" swimtime="00:00:56.36" lane="3" heatid="21010" />
                <RESULT resultid="4693" eventid="23" swimtime="00:03:25.12" lane="2" heatid="23002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:41.40" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1012" birthdate="2011-01-01" gender="F" lastname="Rudolph" firstname="Frieda" license="443387">
              <RESULTS>
                <RESULT resultid="4694" eventid="3" swimtime="00:01:44.07" lane="3" heatid="3006" />
                <RESULT resultid="4695" eventid="10" status="DSQ" swimtime="00:01:30.48" lane="8" heatid="10007" comment="Führte nach verlassen der Rücklage nicht unverzüglich die Wende aus." />
                <RESULT resultid="4696" eventid="14" swimtime="00:03:46.72" lane="8" heatid="14005">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:47.49" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="4697" eventid="19" swimtime="00:00:48.75" lane="8" heatid="19020" />
                <RESULT resultid="4698" eventid="25" swimtime="00:00:40.04" lane="1" heatid="25031" />
                <RESULT resultid="4699" eventid="33" swimtime="00:01:23.57" lane="2" heatid="33011" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1013" birthdate="2007-01-01" gender="F" lastname="Sachs" firstname="Helene" license="344568">
              <RESULTS>
                <RESULT resultid="4700" eventid="3" swimtime="00:01:24.00" lane="5" heatid="3011" />
                <RESULT resultid="4701" eventid="5" swimtime="00:00:33.35" lane="5" heatid="5013" />
                <RESULT resultid="4702" eventid="10" swimtime="00:01:15.36" lane="6" heatid="10016" />
                <RESULT resultid="4703" eventid="14" swimtime="00:03:04.28" lane="5" heatid="14007">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:28.54" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="4704" eventid="33" swimtime="00:01:07.65" lane="4" heatid="33017" />
                <RESULT resultid="4705" eventid="35" swimtime="00:01:24.75" lane="6" heatid="35004" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1014" birthdate="2006-01-01" gender="M" lastname="Bremmers" firstname="Jordi" license="354420">
              <RESULTS>
                <RESULT resultid="4706" eventid="2" swimtime="00:02:25.69" lane="4" heatid="2008">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:08.49" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="4707" eventid="6" swimtime="00:00:27.18" lane="3" heatid="6011" />
                <RESULT resultid="4708" eventid="11" swimtime="00:01:07.92" lane="5" heatid="11012" />
                <RESULT resultid="4709" eventid="13" swimtime="00:00:25.23" lane="4" heatid="13018" />
                <RESULT resultid="4710" eventid="34" swimtime="00:00:57.52" lane="4" heatid="34015" />
                <RESULT resultid="4711" eventid="38" swimtime="00:02:37.93" lane="4" heatid="38005">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:15.15" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1015" birthdate="2015-01-01" gender="M" lastname="Rudolph" firstname="Karl" license="466464">
              <RESULTS>
                <RESULT resultid="4712" eventid="20" swimtime="00:01:10.21" lane="5" heatid="20002" />
                <RESULT resultid="4713" eventid="22" swimtime="00:01:17.81" lane="7" heatid="22003" />
                <RESULT resultid="4714" eventid="26" swimtime="00:00:54.91" lane="6" heatid="26006" />
                <RESULT resultid="4715" eventid="30" swimtime="00:00:51.88" lane="1" heatid="30003" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1016" birthdate="2012-01-01" gender="M" lastname="Winter" firstname="Kevin" license="443384">
              <RESULTS>
                <RESULT resultid="4716" eventid="4" swimtime="00:01:53.26" lane="5" heatid="4003" />
                <RESULT resultid="4717" eventid="11" swimtime="00:01:36.62" lane="2" heatid="11005" />
                <RESULT resultid="4718" eventid="13" swimtime="00:00:37.11" lane="7" heatid="13007" />
                <RESULT resultid="4719" eventid="20" swimtime="00:00:50.32" lane="1" heatid="20013" />
                <RESULT resultid="4720" eventid="24" swimtime="00:03:06.87" lane="7" heatid="24005">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:30.65" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="4721" eventid="34" swimtime="00:01:21.90" lane="6" heatid="34006" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1017" birthdate="2012-01-01" gender="M" lastname="Lindner" firstname="Laurence" license="439928">
              <RESULTS>
                <RESULT resultid="4722" eventid="2" swimtime="00:02:52.41" lane="1" heatid="2007">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:18.92" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="4723" eventid="6" swimtime="00:00:32.80" lane="4" heatid="6008" />
                <RESULT resultid="4724" eventid="11" swimtime="00:01:21.04" lane="2" heatid="11011" />
                <RESULT resultid="4725" eventid="13" swimtime="00:00:32.11" lane="4" heatid="13013" />
                <RESULT resultid="4726" eventid="20" swimtime="00:00:44.63" lane="8" heatid="20018" />
                <RESULT resultid="4727" eventid="24" swimtime="00:02:37.30" lane="8" heatid="24008">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:14.54" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="4728" eventid="26" swimtime="00:00:36.58" lane="4" heatid="26021" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1018" birthdate="2007-01-01" gender="F" lastname="Balkow" firstname="Leonie" license="365625">
              <RESULTS>
                <RESULT resultid="4729" eventid="5" swimtime="00:00:35.09" lane="7" heatid="5012" />
                <RESULT resultid="4730" eventid="12" swimtime="00:00:33.08" lane="4" heatid="12013" />
                <RESULT resultid="4731" eventid="25" swimtime="00:00:37.98" lane="4" heatid="25032" />
                <RESULT resultid="4732" eventid="35" swimtime="00:01:24.20" lane="1" heatid="35004" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1019" birthdate="2011-01-01" gender="M" lastname="Zeretzke" firstname="Linus" license="433193">
              <RESULTS>
                <RESULT resultid="4733" eventid="4" status="DNS" swimtime="00:00:00.00" lane="1" heatid="4009" />
                <RESULT resultid="4734" eventid="13" status="DNS" swimtime="00:00:00.00" lane="5" heatid="13013" />
                <RESULT resultid="4735" eventid="15" status="DNS" swimtime="00:00:00.00" lane="5" heatid="15005" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1020" birthdate="2012-01-01" gender="F" lastname="Wunderlich" firstname="Lotta-Elin" license="436997">
              <RESULTS>
                <RESULT resultid="4736" eventid="1" swimtime="00:02:57.78" lane="5" heatid="1006">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:23.07" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="4737" eventid="5" swimtime="00:00:37.91" lane="4" heatid="5009" />
                <RESULT resultid="4738" eventid="10" swimtime="00:01:25.47" lane="2" heatid="10014" />
                <RESULT resultid="4739" eventid="12" swimtime="00:00:33.86" lane="7" heatid="12013" />
                <RESULT resultid="4740" eventid="23" swimtime="00:02:37.14" lane="7" heatid="23010">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:16.92" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="4741" eventid="25" swimtime="00:00:40.62" lane="3" heatid="25031" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1021" birthdate="2008-01-01" gender="F" lastname="Turczyk" firstname="Lydia" license="349448">
              <RESULTS>
                <RESULT resultid="4742" eventid="5" swimtime="00:00:36.15" lane="4" heatid="5010" />
                <RESULT resultid="4743" eventid="12" swimtime="00:00:33.91" lane="6" heatid="12013" />
                <RESULT resultid="4744" eventid="19" swimtime="00:00:46.66" lane="4" heatid="19020" />
                <RESULT resultid="4745" eventid="25" swimtime="00:00:39.72" lane="6" heatid="25031" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1022" birthdate="2013-01-01" gender="F" lastname="Zeretzke" firstname="Mara" license="455131">
              <RESULTS>
                <RESULT resultid="4746" eventid="3" swimtime="00:01:51.48" lane="4" heatid="3004" />
                <RESULT resultid="4747" eventid="12" swimtime="00:00:40.76" lane="6" heatid="12007" />
                <RESULT resultid="4748" eventid="14" swimtime="00:04:06.30" lane="7" heatid="14003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:58.50" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="4749" eventid="19" swimtime="00:00:49.53" lane="2" heatid="19018" />
                <RESULT resultid="4750" eventid="25" swimtime="00:00:48.72" lane="4" heatid="25018" />
                <RESULT resultid="4751" eventid="31" swimtime="00:01:13.15" lane="3" heatid="31005" />
                <RESULT resultid="4752" eventid="33" swimtime="00:01:37.58" lane="6" heatid="33007" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1023" birthdate="2015-01-01" gender="F" lastname="Künzel" firstname="Marta" license="473898">
              <RESULTS>
                <RESULT resultid="4753" eventid="17" status="DSQ" swimtime="00:01:11.79" lane="8" heatid="17005" comment="Start vor dem Startsignal." />
                <RESULT resultid="4754" eventid="21" status="DSQ" swimtime="00:01:18.93" lane="1" heatid="21004" comment="Das Brett wurde beim Zielanschlag vorn nicht umfasst." />
                <RESULT resultid="4755" eventid="25" swimtime="00:01:04.45" lane="6" heatid="25002" />
                <RESULT resultid="4756" eventid="27" status="DSQ" swimtime="00:01:13.97" lane="3" heatid="27003" comment="Start vor dem Startsignal.&#xA;Wechselbeinschläge nach dem Start." />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1024" birthdate="2013-01-01" gender="M" lastname="Rudert" firstname="Max" license="446075">
              <RESULTS>
                <RESULT resultid="4757" eventid="4" swimtime="00:01:46.55" lane="5" heatid="4006" />
                <RESULT resultid="4758" eventid="11" swimtime="00:01:37.72" lane="7" heatid="11006" />
                <RESULT resultid="4759" eventid="13" swimtime="00:00:37.32" lane="1" heatid="13007" />
                <RESULT resultid="4760" eventid="15" swimtime="00:03:50.49" lane="7" heatid="15004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:51.38" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="4761" eventid="20" swimtime="00:00:47.38" lane="6" heatid="20014" />
                <RESULT resultid="4762" eventid="24" swimtime="00:03:08.75" lane="4" heatid="24005">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:31.21" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="4763" eventid="26" swimtime="00:00:46.09" lane="3" heatid="26017" />
                <RESULT resultid="4764" eventid="34" swimtime="00:01:25.57" lane="7" heatid="34008" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1025" birthdate="2014-01-01" gender="F" lastname="Zwerner" firstname="Nele" license="448863">
              <RESULTS>
                <RESULT resultid="4765" eventid="21" swimtime="00:00:56.20" lane="6" heatid="21012" />
                <RESULT resultid="4766" eventid="25" swimtime="00:00:51.56" lane="1" heatid="25016" />
                <RESULT resultid="4767" eventid="29" swimtime="00:00:43.13" lane="7" heatid="29009" />
                <RESULT resultid="4768" eventid="31" swimtime="00:00:59.40" lane="2" heatid="31006" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1026" birthdate="2014-01-01" gender="M" lastname="Zwerner" firstname="Nils" license="448861">
              <RESULTS>
                <RESULT resultid="4769" eventid="18" swimtime="00:01:07.93" lane="1" heatid="18009" />
                <RESULT resultid="4770" eventid="22" swimtime="00:01:05.04" lane="5" heatid="22007" />
                <RESULT resultid="4771" eventid="26" swimtime="00:00:49.94" lane="8" heatid="26011" />
                <RESULT resultid="4772" eventid="30" swimtime="00:00:42.77" lane="8" heatid="30006" />
                <RESULT resultid="4773" eventid="32" swimtime="00:01:04.40" lane="6" heatid="32003" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1027" birthdate="2013-01-01" gender="M" lastname="Weis" firstname="Simon" license="446189">
              <RESULTS>
                <RESULT resultid="4774" eventid="2" swimtime="00:03:34.92" lane="3" heatid="2003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:41.36" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="4775" eventid="4" swimtime="00:01:57.00" lane="8" heatid="4006" />
                <RESULT resultid="4776" eventid="11" swimtime="00:01:41.12" lane="8" heatid="11005" />
                <RESULT resultid="4777" eventid="13" swimtime="00:00:38.53" lane="7" heatid="13006" />
                <RESULT resultid="4778" eventid="22" swimtime="00:00:59.49" lane="5" heatid="22008" />
                <RESULT resultid="4779" eventid="26" swimtime="00:00:46.47" lane="1" heatid="26016" />
                <RESULT resultid="4780" eventid="34" swimtime="00:01:30.91" lane="2" heatid="34006" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1028" birthdate="2008-01-01" gender="M" lastname="Neumeister" firstname="Til" license="384694">
              <RESULTS>
                <RESULT resultid="4781" eventid="4" swimtime="00:01:19.98" lane="7" heatid="4011" />
                <RESULT resultid="4782" eventid="6" swimtime="00:00:31.34" lane="6" heatid="6010" />
                <RESULT resultid="4783" eventid="13" swimtime="00:00:28.83" lane="1" heatid="13017" />
                <RESULT resultid="4784" eventid="15" swimtime="00:02:58.01" lane="2" heatid="15007">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:23.84" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="4785" eventid="34" swimtime="00:01:05.38" lane="8" heatid="34015" />
                <RESULT resultid="4786" eventid="38" swimtime="00:02:47.31" lane="1" heatid="38005">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:20.29" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1029" birthdate="2015-01-01" gender="M" lastname="Schiller" firstname="Till" license="466462">
              <RESULTS>
                <RESULT resultid="4787" eventid="18" status="DSQ" swimtime="00:01:16.74" lane="8" heatid="18007" comment="Nach dem Start wurde ein Rückenarmzug durchgeführt." />
                <RESULT resultid="4788" eventid="20" swimtime="00:01:08.03" lane="8" heatid="20002" />
                <RESULT resultid="4789" eventid="22" status="DSQ" swimtime="00:01:15.17" lane="2" heatid="22004" comment="2 Brustbeinschläge nach dem Start." />
                <RESULT resultid="4790" eventid="26" swimtime="00:01:01.92" lane="3" heatid="26002" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1030" birthdate="2011-01-01" gender="M" lastname="Schwanke" firstname="Tim" license="423421">
              <RESULTS>
                <RESULT resultid="4791" eventid="11" swimtime="00:01:25.27" lane="1" heatid="11010" />
                <RESULT resultid="4792" eventid="13" swimtime="00:00:30.53" lane="1" heatid="13015" />
                <RESULT resultid="4793" eventid="15" swimtime="00:03:14.87" lane="1" heatid="15006">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:32.86" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="4794" eventid="24" swimtime="00:02:35.45" lane="2" heatid="24008">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:13.06" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="1031" birthdate="2012-01-01" gender="M" lastname="Prager" firstname="Vin-Nino" license="451624">
              <RESULTS>
                <RESULT resultid="4795" eventid="4" swimtime="00:01:41.84" lane="6" heatid="4008" />
                <RESULT resultid="4796" eventid="11" swimtime="00:01:31.86" lane="2" heatid="11008" />
                <RESULT resultid="4797" eventid="15" swimtime="00:03:45.34" lane="2" heatid="15005">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:47.81" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="4798" eventid="22" swimtime="00:00:49.10" lane="3" heatid="22010" />
                <RESULT resultid="4799" eventid="24" swimtime="00:03:05.55" lane="2" heatid="24007">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:26.75" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="4800" eventid="34" swimtime="00:01:20.90" lane="7" heatid="34011" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY number="1" gender="X" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="4677" eventid="16" swimtime="00:02:11.75" lane="5" heatid="16002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:11.94" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1013" number="1" />
                    <RELAYPOSITION athleteid="1028" number="2" />
                    <RELAYPOSITION athleteid="1018" number="3" />
                    <RELAYPOSITION athleteid="1014" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="2" gender="X" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="4678" eventid="7" swimtime="00:02:31.47" lane="1" heatid="7003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:27.17" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1020" number="1" />
                    <RELAYPOSITION athleteid="1031" number="2" />
                    <RELAYPOSITION athleteid="1017" number="3" />
                    <RELAYPOSITION athleteid="1030" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB name="SWV TuR Dresden" nation="GER" region="12" code="3358">
          <ATHLETES>
            <ATHLETE athleteid="721" birthdate="2011-01-01" gender="M" lastname="Bludau" firstname="Tim Bjarte" license="423410">
              <RESULTS>
                <RESULT resultid="3445" eventid="4" swimtime="00:01:24.54" lane="3" heatid="4010" />
                <RESULT resultid="3444" eventid="13" swimtime="00:00:33.17" lane="3" heatid="13009" />
                <RESULT resultid="3443" eventid="15" swimtime="00:03:06.47" lane="4" heatid="15006">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:31.11" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="3442" eventid="20" swimtime="00:00:38.97" lane="6" heatid="20020" />
                <RESULT resultid="3441" eventid="26" swimtime="00:00:38.45" lane="4" heatid="26020" />
                <RESULT resultid="3440" eventid="34" swimtime="00:01:13.70" lane="2" heatid="34010" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="722" birthdate="2015-01-01" gender="F" lastname="Fischer" firstname="Nora" license="465835">
              <RESULTS>
                <RESULT resultid="3449" eventid="19" swimtime="00:00:53.00" lane="6" heatid="19011" />
                <RESULT resultid="3448" eventid="25" swimtime="00:00:50.23" lane="3" heatid="25012" />
                <RESULT resultid="3447" eventid="27" swimtime="00:01:01.06" lane="6" heatid="27010" />
                <RESULT resultid="3446" eventid="29" swimtime="00:00:44.94" lane="3" heatid="29011" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="723" birthdate="2014-01-01" gender="F" lastname="Sillke" firstname="Mina" license="448952">
              <RESULTS>
                <RESULT resultid="3452" eventid="21" swimtime="00:01:04.24" lane="6" heatid="21005" />
                <RESULT resultid="3451" eventid="25" swimtime="00:00:49.36" lane="5" heatid="25014" />
                <RESULT resultid="3450" eventid="29" swimtime="00:00:42.76" lane="6" heatid="29010" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="724" birthdate="2011-01-01" gender="F" lastname="Mauermann" firstname="Mila" license="424568">
              <RESULTS>
                <RESULT resultid="3454" eventid="3" swimtime="00:01:24.04" lane="3" heatid="3011" />
                <RESULT resultid="3453" eventid="10" swimtime="00:01:14.81" lane="3" heatid="10016" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="725" birthdate="2012-01-01" gender="M" lastname="Fischer" firstname="Lennox" license="445086">
              <RESULTS>
                <RESULT resultid="3459" eventid="4" swimtime="00:01:29.69" lane="6" heatid="4009" />
                <RESULT resultid="3458" eventid="15" swimtime="00:03:13.52" lane="2" heatid="15006">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:34.50" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="3457" eventid="20" swimtime="00:00:40.10" lane="8" heatid="20020" />
                <RESULT resultid="3456" eventid="26" swimtime="00:00:37.85" lane="6" heatid="26021" />
                <RESULT resultid="3455" eventid="34" swimtime="00:01:13.86" lane="5" heatid="34011" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="726" birthdate="2009-01-01" gender="F" lastname="Linzmajer" firstname="Lara" license="415694">
              <RESULTS>
                <RESULT resultid="3463" eventid="10" swimtime="00:01:27.93" lane="6" heatid="10010" />
                <RESULT resultid="3462" eventid="12" swimtime="00:00:34.34" lane="6" heatid="12011" />
                <RESULT resultid="3461" eventid="19" swimtime="00:00:46.82" lane="5" heatid="19019" />
                <RESULT resultid="3460" eventid="25" swimtime="00:00:40.34" lane="7" heatid="25029" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="727" birthdate="2006-01-01" gender="M" lastname="Probst" firstname="Kai" license="349820">
              <RESULTS>
                <RESULT resultid="3469" eventid="4" swimtime="00:01:13.00" lane="3" heatid="4011" />
                <RESULT resultid="3468" eventid="6" swimtime="00:00:27.97" lane="6" heatid="6011" />
                <RESULT resultid="3467" eventid="11" swimtime="00:01:07.69" lane="3" heatid="11012" />
                <RESULT resultid="3466" eventid="13" swimtime="00:00:26.24" lane="5" heatid="13018" />
                <RESULT resultid="3465" eventid="20" swimtime="00:00:32.29" lane="4" heatid="20022" />
                <RESULT resultid="3464" eventid="26" swimtime="00:00:30.02" lane="4" heatid="26024" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="728" birthdate="2008-01-01" gender="F" lastname="Opitz" firstname="Juliane" license="366318">
              <RESULTS>
                <RESULT resultid="3474" eventid="5" swimtime="00:00:34.66" lane="7" heatid="5013" />
                <RESULT resultid="3473" eventid="10" swimtime="00:01:21.96" lane="3" heatid="10014" />
                <RESULT resultid="3472" eventid="12" swimtime="00:00:32.58" lane="8" heatid="12017" />
                <RESULT resultid="3471" eventid="19" status="DNS" swimtime="00:00:00.00" lane="1" heatid="19025" />
                <RESULT resultid="3470" eventid="25" status="DNS" swimtime="00:00:00.00" lane="5" heatid="25033" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="729" birthdate="2011-01-01" gender="M" lastname="Riedel" firstname="Fritz" license="423409">
              <RESULTS>
                <RESULT resultid="3477" eventid="6" swimtime="00:00:39.60" lane="5" heatid="6005" />
                <RESULT resultid="3476" eventid="11" swimtime="00:01:37.19" lane="4" heatid="11005" />
                <RESULT resultid="3475" eventid="13" swimtime="00:00:35.86" lane="5" heatid="13007" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="730" birthdate="2014-01-01" gender="F" lastname="Lukoschat" firstname="Franka" license="458407">
              <RESULTS>
                <RESULT resultid="3480" eventid="19" swimtime="00:00:50.86" lane="8" heatid="19015" />
                <RESULT resultid="3479" eventid="25" swimtime="00:00:47.44" lane="2" heatid="25010" />
                <RESULT resultid="3478" eventid="27" swimtime="00:00:59.18" lane="6" heatid="27011" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="731" birthdate="2007-01-01" gender="M" lastname="Dittmar" firstname="Erik" license="364564">
              <RESULTS>
                <RESULT resultid="3488" eventid="2" swimtime="00:02:36.56" lane="2" heatid="2008">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:11.34" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="3487" eventid="6" swimtime="00:00:30.54" lane="1" heatid="6011" />
                <RESULT resultid="3486" eventid="11" swimtime="00:01:11.82" lane="2" heatid="11012" />
                <RESULT resultid="3485" eventid="13" swimtime="00:00:28.57" lane="7" heatid="13017" />
                <RESULT resultid="3484" eventid="20" swimtime="00:00:36.80" lane="1" heatid="20022" />
                <RESULT resultid="3483" eventid="26" swimtime="00:00:32.51" lane="2" heatid="26024" />
                <RESULT resultid="3482" eventid="34" swimtime="00:01:02.72" lane="7" heatid="34015" />
                <RESULT resultid="3481" eventid="38" status="DNS" swimtime="00:00:00.00" lane="6" heatid="38005" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="732" birthdate="2009-01-01" gender="M" lastname="Mätzold" firstname="Collin" license="371200">
              <RESULTS>
                <RESULT resultid="3491" eventid="20" swimtime="00:00:42.55" lane="7" heatid="20018" />
                <RESULT resultid="3490" eventid="24" swimtime="00:02:54.22" lane="4" heatid="24006">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:19.52" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="3489" eventid="26" swimtime="00:00:37.54" lane="3" heatid="26021" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="733" birthdate="2013-01-01" gender="F" lastname="Mätzold" firstname="Chiara" license="448443">
              <RESULTS>
                <RESULT resultid="3494" eventid="17" swimtime="00:01:07.25" lane="6" heatid="17010" />
                <RESULT resultid="3493" eventid="21" swimtime="00:01:08.77" lane="7" heatid="21009" />
                <RESULT resultid="3492" eventid="25" swimtime="00:00:48.63" lane="2" heatid="25013" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="734" birthdate="2013-01-01" gender="M" lastname="Mätzold" firstname="Chris" license="448442">
              <RESULTS>
                <RESULT resultid="3497" eventid="20" swimtime="00:00:54.44" lane="8" heatid="20009" />
                <RESULT resultid="3496" eventid="26" swimtime="00:01:01.79" lane="7" heatid="26004" />
                <RESULT resultid="3495" eventid="28" swimtime="00:01:03.36" lane="2" heatid="28006" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY number="1" gender="X" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="3498" eventid="7" swimtime="00:02:23.12" lane="7" heatid="7003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:16.88" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="725" number="1" />
                    <RELAYPOSITION athleteid="721" number="2" />
                    <RELAYPOSITION athleteid="724" number="3" />
                    <RELAYPOSITION athleteid="729" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" gender="X" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="3499" eventid="16" swimtime="00:02:10.42" lane="2" heatid="16002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:04.31" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="731" number="1" />
                    <RELAYPOSITION athleteid="727" number="2" />
                    <RELAYPOSITION athleteid="728" number="3" />
                    <RELAYPOSITION athleteid="732" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB name="Tauchclub NEMO Plauen e.V." nation="GER" region="20" code="0">
          <ATHLETES>
            <ATHLETE athleteid="103" birthdate="2012-01-01" gender="M" lastname="Ngo" firstname="Charlie James" license="0">
              <RESULTS>
                <RESULT resultid="565" eventid="40" swimtime="00:03:12.02" lane="1" heatid="40002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:38.71" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="566" eventid="42" status="DSQ" swimtime="00:00:22.37" lane="5" heatid="42001" comment="Gesicht aus dem Wasser." />
                <RESULT resultid="567" eventid="46" swimtime="00:01:25.20" lane="1" heatid="46002" />
                <RESULT resultid="568" eventid="50" swimtime="00:00:34.26" lane="6" heatid="50002" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="104" birthdate="2013-01-01" gender="M" lastname="Hertel" firstname="Etienne" license="0">
              <RESULTS>
                <RESULT resultid="569" eventid="40" swimtime="00:02:53.81" lane="4" heatid="40001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:21.52" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="570" eventid="42" swimtime="00:00:19.54" lane="4" heatid="42001" />
                <RESULT resultid="571" eventid="46" swimtime="00:01:24.52" lane="2" heatid="46001" />
                <RESULT resultid="572" eventid="50" swimtime="00:00:35.90" lane="4" heatid="50001" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="105" birthdate="2011-01-01" gender="F" lastname="Köhler" firstname="Josephine" license="0">
              <RESULTS>
                <RESULT resultid="573" eventid="39" swimtime="00:03:24.94" lane="3" heatid="39001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:31.30" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="574" eventid="45" swimtime="00:01:34.64" lane="2" heatid="45002" />
                <RESULT resultid="575" eventid="49" swimtime="00:00:40.34" lane="4" heatid="49001" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="106" birthdate="2010-01-01" gender="F" lastname="Dawert" firstname="Klara" license="0">
              <RESULTS>
                <RESULT resultid="576" eventid="41" swimtime="00:00:16.74" lane="6" heatid="41001" />
                <RESULT resultid="577" eventid="45" swimtime="00:01:12.33" lane="6" heatid="45004" />
                <RESULT resultid="578" eventid="49" swimtime="00:00:33.34" lane="1" heatid="49003" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="107" birthdate="2013-01-01" gender="F" lastname="Küthemann" firstname="Lina" license="0">
              <RESULTS>
                <RESULT resultid="579" eventid="39" swimtime="00:02:45.57" lane="5" heatid="39001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:19.81" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="580" eventid="41" swimtime="00:00:15.71" lane="3" heatid="41001" />
                <RESULT resultid="581" eventid="45" swimtime="00:01:13.55" lane="8" heatid="45003" />
                <RESULT resultid="582" eventid="49" swimtime="00:00:32.97" lane="6" heatid="49002" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="108" birthdate="2008-01-01" gender="F" lastname="Weller" firstname="Maren" license="0">
              <RESULTS>
                <RESULT resultid="583" eventid="39" swimtime="00:02:25.14" lane="6" heatid="39002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:08.53" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="584" eventid="41" swimtime="00:00:15.81" lane="3" heatid="41003" />
                <RESULT resultid="585" eventid="45" swimtime="00:01:01.59" lane="1" heatid="45006" />
                <RESULT resultid="586" eventid="49" swimtime="00:00:27.80" lane="5" heatid="49004" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="109" birthdate="2014-01-01" gender="M" lastname="Michalke" firstname="Max-Leon" license="0">
              <RESULTS>
                <RESULT resultid="587" eventid="40" swimtime="00:03:00.66" lane="7" heatid="40002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:27.88" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="588" eventid="44" swimtime="00:00:18.38" lane="4" heatid="44001" />
                <RESULT resultid="589" eventid="46" swimtime="00:01:27.33" lane="8" heatid="46002" />
                <RESULT resultid="590" eventid="50" swimtime="00:00:37.24" lane="7" heatid="50002" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="110" birthdate="2013-01-01" gender="M" lastname="Hartmann" firstname="Paul" license="0">
              <RESULTS>
                <RESULT resultid="591" eventid="40" swimtime="00:02:26.86" lane="6" heatid="40002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:17.64" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="592" eventid="42" swimtime="00:00:16.07" lane="2" heatid="42002" />
                <RESULT resultid="593" eventid="46" swimtime="00:01:19.03" lane="5" heatid="46002" />
                <RESULT resultid="594" eventid="50" swimtime="00:00:32.72" lane="1" heatid="50003" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="111" birthdate="2008-01-01" gender="F" lastname="Steinert" firstname="Sara-Marie" license="0">
              <RESULTS>
                <RESULT resultid="595" eventid="39" swimtime="00:03:40.42" lane="6" heatid="39001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:43.83" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="596" eventid="41" status="DSQ" swimtime="00:00:40.25" lane="2" heatid="41001" comment="Aufgegeben nach 10 Meter." />
                <RESULT resultid="597" eventid="45" swimtime="00:01:43.16" lane="4" heatid="45001" />
                <RESULT resultid="598" eventid="49" swimtime="00:00:42.36" lane="5" heatid="49001" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="112" birthdate="2010-01-01" gender="F" lastname="Martin" firstname="Theresa" license="0">
              <RESULTS>
                <RESULT resultid="599" eventid="39" swimtime="00:02:29.03" lane="8" heatid="39003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:08.10" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="600" eventid="41" swimtime="00:00:15.68" lane="2" heatid="41003" />
                <RESULT resultid="601" eventid="45" swimtime="00:01:04.39" lane="2" heatid="45005" />
                <RESULT resultid="602" eventid="49" swimtime="00:00:28.86" lane="7" heatid="49004" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="113" birthdate="2007-01-01" gender="M" lastname="Kaden" firstname="Tim" license="0">
              <RESULTS>
                <RESULT resultid="603" eventid="40" swimtime="00:02:30.71" lane="3" heatid="40002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:11.66" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="604" eventid="46" swimtime="00:01:03.56" lane="7" heatid="46003" />
                <RESULT resultid="605" eventid="50" swimtime="00:00:27.78" lane="3" heatid="50003" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="114" birthdate="2013-01-01" gender="M" lastname="Kad" firstname="Vincent" license="0">
              <RESULTS>
                <RESULT resultid="606" eventid="40" swimtime="00:03:00.12" lane="8" heatid="40002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:28.63" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="607" eventid="42" swimtime="00:00:20.50" lane="3" heatid="42001" />
                <RESULT resultid="608" eventid="46" swimtime="00:01:23.37" lane="5" heatid="46001" />
                <RESULT resultid="609" eventid="50" swimtime="00:00:36.90" lane="8" heatid="50002" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="TC Delitzsch" nation="GER" region="20" code="0">
          <ATHLETES>
            <ATHLETE athleteid="445" birthdate="2011-01-01" gender="M" lastname="Becker" firstname="Pepe Milan" license="0">
              <RESULTS>
                <RESULT resultid="2148" eventid="40" swimtime="00:02:11.34" lane="5" heatid="40002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:05.34" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="2147" eventid="42" swimtime="00:00:13.57" lane="6" heatid="42003" />
                <RESULT resultid="2146" eventid="46" swimtime="00:00:59.71" lane="6" heatid="46003" />
                <RESULT resultid="2145" eventid="48" swimtime="00:00:40.80" lane="1" heatid="48001" />
                <RESULT resultid="2144" eventid="50" swimtime="00:00:25.75" lane="5" heatid="50003" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="446" birthdate="2011-01-01" gender="F" lastname="Schönherr" firstname="Nina" license="0">
              <RESULTS>
                <RESULT resultid="2153" eventid="39" swimtime="00:02:16.57" lane="6" heatid="39003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:03.57" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="2152" eventid="41" swimtime="00:00:14.58" lane="6" heatid="41005" />
                <RESULT resultid="2151" eventid="45" swimtime="00:00:59.55" lane="3" heatid="45006" />
                <RESULT resultid="2150" eventid="47" swimtime="00:00:36.33" lane="5" heatid="47001" />
                <RESULT resultid="2149" eventid="49" swimtime="00:00:26.52" lane="6" heatid="49005" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="USV TU Dresden e.V." nation="GER" region="12" code="3410">
          <ATHLETES>
            <ATHLETE athleteid="385" birthdate="2015-01-01" gender="M" lastname="Hebold" firstname="Toni" license="453990">
              <RESULTS>
                <RESULT resultid="1886" eventid="18" swimtime="00:01:19.84" lane="3" heatid="18005" />
                <RESULT resultid="1885" eventid="22" swimtime="00:01:19.39" lane="8" heatid="22003" />
                <RESULT resultid="1884" eventid="26" swimtime="00:00:59.76" lane="7" heatid="26002" />
                <RESULT resultid="1883" eventid="30" swimtime="00:01:03.29" lane="8" heatid="30002" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="386" birthdate="2010-01-01" gender="M" lastname="Kobsch" firstname="Tim-Ruben" license="456815">
              <RESULTS>
                <RESULT resultid="1890" eventid="20" swimtime="00:00:51.19" lane="2" heatid="20010" />
                <RESULT resultid="1889" eventid="24" swimtime="00:03:14.91" lane="3" heatid="24003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:35.92" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1888" eventid="26" swimtime="00:00:48.78" lane="6" heatid="26013" />
                <RESULT resultid="1887" eventid="34" swimtime="00:01:27.44" lane="6" heatid="34004" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="387" birthdate="2012-01-01" gender="F" lastname="Einbock" firstname="Theresa" license="445207">
              <RESULTS>
                <RESULT resultid="1895" eventid="12" swimtime="00:00:35.68" lane="5" heatid="12007" />
                <RESULT resultid="1894" eventid="14" swimtime="00:03:22.34" lane="5" heatid="14005">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:37.41" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1893" eventid="19" swimtime="00:00:41.74" lane="3" heatid="19023" />
                <RESULT resultid="1892" eventid="23" swimtime="00:03:11.85" lane="1" heatid="23003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:31.46" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1891" eventid="25" swimtime="00:00:44.97" lane="4" heatid="25022" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="388" birthdate="2015-01-01" gender="M" lastname="Grams" firstname="Sascha" license="471326">
              <RESULTS>
                <RESULT resultid="1899" eventid="18" swimtime="00:01:14.81" lane="4" heatid="18003" />
                <RESULT resultid="1898" eventid="20" swimtime="00:00:58.32" lane="2" heatid="20005" />
                <RESULT resultid="1897" eventid="26" swimtime="00:01:00.14" lane="6" heatid="26002" />
                <RESULT resultid="1896" eventid="28" swimtime="00:01:08.69" lane="6" heatid="28003" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="389" birthdate="2015-01-01" gender="F" lastname="Küng" firstname="Ronja" license="472898">
              <RESULTS>
                <RESULT resultid="1904" eventid="17" status="DSQ" swimtime="00:01:23.49" lane="2" heatid="17003" comment="Rückenarmbewegung nach dem Start." />
                <RESULT resultid="1903" eventid="19" swimtime="00:01:00.44" lane="5" heatid="19001" />
                <RESULT resultid="1902" eventid="21" swimtime="00:01:11.49" lane="2" heatid="21003" />
                <RESULT resultid="1901" eventid="25" swimtime="00:01:10.69" lane="4" heatid="25002" />
                <RESULT resultid="1900" eventid="27" swimtime="00:01:11.02" lane="6" heatid="27003" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="390" birthdate="2014-01-01" gender="F" lastname="Plietker" firstname="Ria Johanna" license="448836">
              <RESULTS>
                <RESULT resultid="1909" eventid="17" swimtime="00:01:06.30" lane="2" heatid="17008" />
                <RESULT resultid="1908" eventid="19" swimtime="00:00:53.32" lane="8" heatid="19013" />
                <RESULT resultid="1907" eventid="25" swimtime="00:00:50.52" lane="7" heatid="25009" />
                <RESULT resultid="1906" eventid="29" swimtime="00:00:44.34" lane="8" heatid="29009" />
                <RESULT resultid="1905" eventid="33" swimtime="00:01:38.37" lane="3" heatid="33003" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="391" birthdate="2007-01-01" gender="F" lastname="Schmidt" firstname="Paula" license="376891">
              <RESULTS>
                <RESULT resultid="1912" eventid="1" swimtime="00:03:23.89" lane="3" heatid="1003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:36.46" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1911" eventid="10" swimtime="00:01:25.12" lane="2" heatid="10012" />
                <RESULT resultid="1910" eventid="12" swimtime="00:00:33.28" lane="4" heatid="12011" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="392" birthdate="2010-01-01" gender="F" lastname="Rülker" firstname="Nina" license="437636">
              <RESULTS>
                <RESULT resultid="1915" eventid="23" swimtime="00:02:47.52" lane="7" heatid="23007">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:20.74" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1914" eventid="33" swimtime="00:01:15.65" lane="1" heatid="33014" />
                <RESULT resultid="1913" eventid="37" swimtime="00:03:21.59" lane="7" heatid="37002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:38.48" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="393" birthdate="2013-01-01" gender="F" lastname="Kern" firstname="Nieke" license="447949">
              <RESULTS>
                <RESULT resultid="1921" eventid="10" swimtime="00:01:33.87" lane="4" heatid="10009" />
                <RESULT resultid="1920" eventid="12" swimtime="00:00:40.25" lane="8" heatid="12007" />
                <RESULT resultid="1919" eventid="17" swimtime="00:00:52.25" lane="1" heatid="17015" />
                <RESULT resultid="1918" eventid="25" swimtime="00:00:42.04" lane="8" heatid="25027" />
                <RESULT resultid="1917" eventid="33" swimtime="00:01:33.96" lane="7" heatid="33008" />
                <RESULT resultid="1916" eventid="37" swimtime="00:03:26.22" lane="7" heatid="37003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:39.93" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="394" birthdate="2009-01-01" gender="F" lastname="Tasarz" firstname="Nida" license="460651">
              <RESULTS>
                <RESULT resultid="1924" eventid="23" swimtime="00:03:04.48" lane="2" heatid="23005">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:25.50" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1923" eventid="25" swimtime="00:00:43.54" lane="1" heatid="25025" />
                <RESULT resultid="1922" eventid="33" swimtime="00:01:26.09" lane="5" heatid="33008" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="395" birthdate="2015-01-01" gender="F" lastname="Mühlenberg" firstname="Nele" license="471480">
              <RESULTS>
                <RESULT resultid="1928" eventid="17" swimtime="00:01:15.71" lane="4" heatid="17001" />
                <RESULT resultid="1927" eventid="19" swimtime="00:01:08.86" lane="8" heatid="19002" />
                <RESULT resultid="1926" eventid="25" swimtime="00:01:14.51" lane="7" heatid="25002" />
                <RESULT resultid="1925" eventid="27" swimtime="00:01:16.50" lane="8" heatid="27003" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="396" birthdate="2010-01-01" gender="M" lastname="Jacob" firstname="Moritz" license="410639">
              <RESULTS>
                <RESULT resultid="1934" eventid="2" swimtime="00:03:21.18" lane="8" heatid="2003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:36.63" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1933" eventid="11" swimtime="00:01:29.42" lane="4" heatid="11008" />
                <RESULT resultid="1932" eventid="13" swimtime="00:00:35.99" lane="5" heatid="13005" />
                <RESULT resultid="1931" eventid="20" swimtime="00:00:48.26" lane="8" heatid="20010" />
                <RESULT resultid="1930" eventid="26" swimtime="00:00:40.82" lane="4" heatid="26016" />
                <RESULT resultid="1929" eventid="38" swimtime="00:03:10.31" lane="5" heatid="38003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:34.82" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="397" birthdate="2011-01-01" gender="M" lastname="Schwarzer" firstname="Max" license="437639">
              <RESULTS>
                <RESULT resultid="1938" eventid="11" swimtime="00:01:27.22" lane="6" heatid="11009" />
                <RESULT resultid="1937" eventid="13" swimtime="00:00:34.58" lane="8" heatid="13010" />
                <RESULT resultid="1936" eventid="34" swimtime="00:01:19.08" lane="2" heatid="34009" />
                <RESULT resultid="1935" eventid="38" swimtime="00:03:06.99" lane="6" heatid="38003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:30.61" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="398" birthdate="2014-01-01" gender="F" lastname="Krusch" firstname="Mathilda" license="459676">
              <RESULTS>
                <RESULT resultid="1943" eventid="17" swimtime="00:01:15.77" lane="7" heatid="17005" />
                <RESULT resultid="1942" eventid="19" swimtime="00:01:02.89" lane="5" heatid="19005" />
                <RESULT resultid="1941" eventid="25" swimtime="00:01:03.19" lane="8" heatid="25003" />
                <RESULT resultid="1940" eventid="27" swimtime="00:01:11.26" lane="5" heatid="27003" />
                <RESULT resultid="1939" eventid="29" swimtime="00:01:03.27" lane="1" heatid="29002" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="399" birthdate="2010-01-01" gender="F" lastname="Birn" firstname="Marie Luise" license="426670">
              <RESULTS>
                <RESULT resultid="1948" eventid="1" swimtime="00:03:07.10" lane="2" heatid="1002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:26.60" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1947" eventid="10" swimtime="00:01:30.86" lane="3" heatid="10006" />
                <RESULT resultid="1946" eventid="12" swimtime="00:00:34.56" lane="3" heatid="12010" />
                <RESULT resultid="1945" eventid="23" swimtime="00:02:44.66" lane="8" heatid="23004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:20.48" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1944" eventid="33" swimtime="00:01:14.11" lane="1" heatid="33011" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="400" birthdate="2012-01-01" gender="F" lastname="Schumann" firstname="Margot" license="437638">
              <RESULTS>
                <RESULT resultid="1953" eventid="12" swimtime="00:00:39.16" lane="2" heatid="12005" />
                <RESULT resultid="1952" eventid="14" swimtime="00:03:34.91" lane="3" heatid="14004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:44.43" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1951" eventid="19" swimtime="00:00:44.11" lane="4" heatid="19021" />
                <RESULT resultid="1950" eventid="23" swimtime="00:03:20.35" lane="6" heatid="23001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:36.50" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1949" eventid="25" swimtime="00:00:43.28" lane="2" heatid="25022" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="401" birthdate="2012-01-01" gender="F" lastname="Dittel" firstname="Magdalena" license="437623">
              <RESULTS>
                <RESULT resultid="1957" eventid="5" swimtime="00:00:36.85" lane="8" heatid="5011" />
                <RESULT resultid="1956" eventid="14" swimtime="00:03:38.42" lane="5" heatid="14001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:46.27" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1955" eventid="23" swimtime="00:02:36.22" lane="6" heatid="23010">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:16.00" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1954" eventid="35" swimtime="00:01:29.95" lane="2" heatid="35003" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="402" birthdate="2011-01-01" gender="M" lastname="Ranft" firstname="Lukas" license="426681">
              <RESULTS>
                <RESULT resultid="1960" eventid="2" status="WDR" swimtime="00:00:00.00" lane="5" heatid="2002" />
                <RESULT resultid="1959" eventid="11" status="WDR" swimtime="00:00:00.00" lane="4" heatid="11007" />
                <RESULT resultid="1958" eventid="13" status="WDR" swimtime="00:00:00.00" lane="8" heatid="13012" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="403" birthdate="2011-01-01" gender="M" lastname="Langner" firstname="Lukas" license="426678">
              <RESULTS>
                <RESULT resultid="1962" eventid="4" swimtime="00:01:29.46" lane="2" heatid="4009" />
                <RESULT resultid="1961" eventid="9" swimtime="00:02:50.43" lane="6" heatid="9001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:19.41" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="404" birthdate="2013-01-01" gender="F" lastname="Prager" firstname="Luise" license="451488">
              <RESULTS>
                <RESULT resultid="1966" eventid="19" swimtime="00:01:03.08" lane="7" heatid="19005" />
                <RESULT resultid="1965" eventid="21" swimtime="00:01:20.69" lane="3" heatid="21002" />
                <RESULT resultid="1964" eventid="25" swimtime="00:01:01.27" lane="6" heatid="25003" />
                <RESULT resultid="1963" eventid="33" swimtime="00:02:15.63" lane="4" heatid="33001" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="405" birthdate="2014-01-01" gender="M" lastname="Sacher" firstname="Louis" license="459819">
              <RESULTS>
                <RESULT resultid="1971" eventid="18" swimtime="00:01:05.34" lane="3" heatid="18009" />
                <RESULT resultid="1970" eventid="20" swimtime="00:00:57.40" lane="5" heatid="20006" />
                <RESULT resultid="1969" eventid="26" swimtime="00:00:49.64" lane="1" heatid="26011" />
                <RESULT resultid="1968" eventid="30" swimtime="00:00:44.28" lane="7" heatid="30007" />
                <RESULT resultid="1967" eventid="34" swimtime="00:01:41.59" lane="6" heatid="34002" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="406" birthdate="2015-01-01" gender="F" lastname="Grumbt" firstname="Lisa" license="468359">
              <RESULTS>
                <RESULT resultid="1976" eventid="17" swimtime="00:01:09.50" lane="6" heatid="17014" />
                <RESULT resultid="1975" eventid="19" swimtime="00:01:06.43" lane="1" heatid="19003" />
                <RESULT resultid="1974" eventid="21" swimtime="00:01:02.93" lane="5" heatid="21010" />
                <RESULT resultid="1973" eventid="25" swimtime="00:00:54.67" lane="8" heatid="25009" />
                <RESULT resultid="1972" eventid="29" swimtime="00:00:51.98" lane="7" heatid="29006" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="407" birthdate="2015-01-01" gender="F" lastname="Pouva" firstname="Lilli" license="463785">
              <RESULTS>
                <RESULT resultid="1981" eventid="17" swimtime="00:01:13.13" lane="2" heatid="17009" />
                <RESULT resultid="1980" eventid="19" swimtime="00:01:03.28" lane="5" heatid="19003" />
                <RESULT resultid="1979" eventid="25" swimtime="00:00:56.41" lane="5" heatid="25006" />
                <RESULT resultid="1978" eventid="27" swimtime="00:01:19.18" lane="5" heatid="27004" />
                <RESULT resultid="1977" eventid="29" swimtime="00:00:56.48" lane="8" heatid="29004" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="408" birthdate="2010-01-01" gender="M" lastname="Tkachenko" firstname="Leonard" license="410656">
              <RESULTS>
                <RESULT resultid="1984" eventid="24" swimtime="00:03:00.99" lane="4" heatid="24004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:26.19" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1983" eventid="34" swimtime="00:01:22.76" lane="5" heatid="34008" />
                <RESULT resultid="1982" eventid="38" swimtime="00:03:23.37" lane="2" heatid="38002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:40.46" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="409" birthdate="2011-01-01" gender="F" lastname="Maihold" firstname="Lea-Sophie" license="437630">
              <RESULTS>
                <RESULT resultid="1989" eventid="12" swimtime="00:00:33.92" lane="1" heatid="12010" />
                <RESULT resultid="1988" eventid="14" swimtime="00:03:37.30" lane="1" heatid="14002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:45.09" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1987" eventid="19" swimtime="00:00:46.35" lane="3" heatid="19019" />
                <RESULT resultid="1986" eventid="23" swimtime="00:03:04.66" lane="1" heatid="23004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:27.03" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1985" eventid="37" swimtime="00:03:11.96" lane="8" heatid="37002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:34.94" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="410" birthdate="2012-01-01" gender="F" lastname="Eisert" firstname="Lea" license="437624">
              <RESULTS>
                <RESULT resultid="1994" eventid="10" swimtime="00:01:27.38" lane="3" heatid="10012" />
                <RESULT resultid="1993" eventid="12" swimtime="00:00:33.60" lane="7" heatid="12014" />
                <RESULT resultid="1992" eventid="23" swimtime="00:02:51.50" lane="1" heatid="23006">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:24.13" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1991" eventid="25" swimtime="00:00:39.83" lane="4" heatid="25031" />
                <RESULT resultid="1990" eventid="37" swimtime="00:03:05.41" lane="1" heatid="37005">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:31.91" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="411" birthdate="2013-01-01" gender="F" lastname="Neubauer" firstname="Laila" license="447951">
              <RESULTS>
                <RESULT resultid="1998" eventid="19" swimtime="00:00:51.53" lane="8" heatid="19012" />
                <RESULT resultid="1997" eventid="25" swimtime="00:00:52.24" lane="7" heatid="25014" />
                <RESULT resultid="1996" eventid="27" swimtime="00:01:06.39" lane="3" heatid="27005" />
                <RESULT resultid="1995" eventid="33" swimtime="00:01:48.74" lane="8" heatid="33003" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="412" birthdate="2014-01-01" gender="M" lastname="Labuschke" firstname="Konstantin" license="451949">
              <RESULTS>
                <RESULT resultid="2003" eventid="18" swimtime="00:00:59.79" lane="2" heatid="18010" />
                <RESULT resultid="2002" eventid="22" swimtime="00:00:55.87" lane="1" heatid="22010" />
                <RESULT resultid="2001" eventid="26" swimtime="00:00:49.45" lane="4" heatid="26008" />
                <RESULT resultid="2000" eventid="30" swimtime="00:00:44.75" lane="1" heatid="30006" />
                <RESULT resultid="1999" eventid="32" swimtime="00:01:06.41" lane="4" heatid="32002" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="413" birthdate="2012-01-01" gender="M" lastname="Kurlykov" firstname="Kirill" license="437629">
              <RESULTS>
                <RESULT resultid="2009" eventid="11" swimtime="00:01:23.80" lane="2" heatid="11009" />
                <RESULT resultid="2008" eventid="15" swimtime="00:03:27.21" lane="1" heatid="15005">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:40.20" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="2007" eventid="20" swimtime="00:00:44.39" lane="4" heatid="20017" />
                <RESULT resultid="2006" eventid="28" swimtime="00:00:55.65" lane="6" heatid="28007" />
                <RESULT resultid="2005" eventid="34" swimtime="00:01:14.65" lane="4" heatid="34011" />
                <RESULT resultid="2004" eventid="38" swimtime="00:03:04.01" lane="8" heatid="38003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:31.90" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="414" birthdate="2008-01-01" gender="F" lastname="Grammlich" firstname="Katharina" license="380800">
              <RESULTS>
                <RESULT resultid="2012" eventid="10" swimtime="00:01:08.50" lane="4" heatid="10016" />
                <RESULT resultid="2011" eventid="25" swimtime="00:00:31.34" lane="4" heatid="25034" />
                <RESULT resultid="2010" eventid="37" swimtime="00:02:29.04" lane="4" heatid="37007">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:13.25" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="415" birthdate="2014-01-01" gender="F" lastname="Six" firstname="Juli" license="459728">
              <RESULTS>
                <RESULT resultid="2017" eventid="17" swimtime="00:01:04.23" lane="2" heatid="17010" />
                <RESULT resultid="2016" eventid="21" swimtime="00:01:11.69" lane="6" heatid="21006" />
                <RESULT resultid="2015" eventid="25" swimtime="00:00:50.01" lane="8" heatid="25017" />
                <RESULT resultid="2014" eventid="29" swimtime="00:00:50.05" lane="5" heatid="29007" />
                <RESULT resultid="2013" eventid="33" swimtime="00:01:52.13" lane="6" heatid="33002" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="416" birthdate="2014-01-01" gender="M" lastname="Ranft" firstname="Jonas" license="451486">
              <RESULTS>
                <RESULT resultid="2022" eventid="18" swimtime="00:01:18.40" lane="4" heatid="18002" />
                <RESULT resultid="2021" eventid="20" swimtime="00:01:03.22" lane="2" heatid="20003" />
                <RESULT resultid="2020" eventid="22" swimtime="00:01:25.70" lane="3" heatid="22001" />
                <RESULT resultid="2019" eventid="28" swimtime="00:01:10.49" lane="7" heatid="28002" />
                <RESULT resultid="2018" eventid="30" swimtime="00:01:00.88" lane="4" heatid="30001" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="417" birthdate="2010-01-01" gender="M" lastname="Höhne" firstname="Janek" license="410637">
              <RESULTS>
                <RESULT resultid="2025" eventid="2" swimtime="00:03:19.78" lane="8" heatid="2004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:39.30" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="2024" eventid="11" swimtime="00:01:37.75" lane="8" heatid="11008" />
                <RESULT resultid="2023" eventid="13" swimtime="00:00:36.79" lane="2" heatid="13010" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="418" birthdate="2015-01-01" gender="M" lastname="Litta" firstname="Henrik" license="463806">
              <RESULTS>
                <RESULT resultid="2030" eventid="20" swimtime="00:00:58.42" lane="6" heatid="20008" />
                <RESULT resultid="2029" eventid="22" status="DSQ" swimtime="00:01:06.47" lane="2" heatid="22007" comment="Start vor dem Startsignal." />
                <RESULT resultid="2028" eventid="26" swimtime="00:00:51.56" lane="5" heatid="26007" />
                <RESULT resultid="2027" eventid="28" swimtime="00:01:12.97" lane="4" heatid="28004" />
                <RESULT resultid="2026" eventid="30" swimtime="00:00:49.78" lane="6" heatid="30005" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="419" birthdate="2011-01-01" gender="F" lastname="Rex" firstname="Henriette" license="426682">
              <RESULTS>
                <RESULT resultid="2033" eventid="23" swimtime="00:02:52.32" lane="7" heatid="23008">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:21.57" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="2032" eventid="33" swimtime="00:01:17.88" lane="4" heatid="33012" />
                <RESULT resultid="2031" eventid="37" swimtime="00:03:11.98" lane="3" heatid="37003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:35.01" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="420" birthdate="2013-01-01" gender="M" lastname="Lutter" firstname="Henning" license="445208">
              <RESULTS>
                <RESULT resultid="2037" eventid="20" swimtime="00:00:57.13" lane="7" heatid="20006" />
                <RESULT resultid="2036" eventid="22" swimtime="00:01:06.43" lane="6" heatid="22007" />
                <RESULT resultid="2035" eventid="26" swimtime="00:00:49.87" lane="2" heatid="26010" />
                <RESULT resultid="2034" eventid="34" swimtime="00:01:33.35" lane="2" heatid="34003" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="421" birthdate="2015-01-01" gender="F" lastname="Westphal" firstname="Helen" license="464958">
              <RESULTS>
                <RESULT resultid="2041" eventid="17" status="DNS" swimtime="00:00:00.00" lane="7" heatid="17002" />
                <RESULT resultid="2040" eventid="19" status="DNS" swimtime="00:00:00.00" lane="3" heatid="19001" />
                <RESULT resultid="2039" eventid="25" status="DNS" swimtime="00:00:00.00" lane="5" heatid="25002" />
                <RESULT resultid="2038" eventid="27" status="DNS" swimtime="00:00:00.00" lane="1" heatid="27003" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="422" birthdate="2007-01-01" gender="F" lastname="Kiontke" firstname="Franziska" license="364576">
              <RESULTS>
                <RESULT resultid="2044" eventid="23" status="WDR" swimtime="00:00:00.00" lane="8" heatid="23007" />
                <RESULT resultid="2043" eventid="33" status="WDR" swimtime="00:00:00.00" lane="8" heatid="33015" />
                <RESULT resultid="2042" eventid="37" status="WDR" swimtime="00:00:00.00" lane="7" heatid="37004" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="423" birthdate="2010-01-01" gender="M" lastname="Tröger" firstname="Florian" license="426687">
              <RESULTS>
                <RESULT resultid="2048" eventid="20" swimtime="00:00:45.64" lane="7" heatid="20013" />
                <RESULT resultid="2047" eventid="24" swimtime="00:03:14.19" lane="5" heatid="24003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:28.92" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="2046" eventid="26" swimtime="00:00:43.61" lane="6" heatid="26014" />
                <RESULT resultid="2045" eventid="34" swimtime="00:01:25.61" lane="4" heatid="34004" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="424" birthdate="2014-01-01" gender="M" lastname="Scholz" firstname="Ferdinand" license="456406">
              <RESULTS>
                <RESULT resultid="2053" eventid="18" swimtime="00:01:08.57" lane="8" heatid="18005" />
                <RESULT resultid="2052" eventid="20" swimtime="00:01:03.56" lane="7" heatid="20003" />
                <RESULT resultid="2051" eventid="22" swimtime="00:01:08.15" lane="7" heatid="22006" />
                <RESULT resultid="2050" eventid="26" swimtime="00:00:56.32" lane="6" heatid="26004" />
                <RESULT resultid="2049" eventid="30" swimtime="00:00:55.32" lane="6" heatid="30002" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="425" birthdate="2014-01-01" gender="M" lastname="Müller" firstname="Felix" license="447956">
              <RESULTS>
                <RESULT resultid="2058" eventid="20" swimtime="00:00:52.56" lane="5" heatid="20011" />
                <RESULT resultid="2057" eventid="22" swimtime="00:00:54.26" lane="3" heatid="22008" />
                <RESULT resultid="2056" eventid="26" swimtime="00:00:44.81" lane="7" heatid="26016" />
                <RESULT resultid="2055" eventid="30" swimtime="00:00:37.77" lane="4" heatid="30008" />
                <RESULT resultid="2054" eventid="34" swimtime="00:01:29.42" lane="4" heatid="34003" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="426" birthdate="2011-01-01" gender="F" lastname="Schumann" firstname="Ella" license="426684">
              <RESULTS>
                <RESULT resultid="2064" eventid="1" swimtime="00:03:15.61" lane="7" heatid="1003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:30.97" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="2063" eventid="10" swimtime="00:01:30.94" lane="1" heatid="10009" />
                <RESULT resultid="2062" eventid="12" swimtime="00:00:35.29" lane="1" heatid="12009" />
                <RESULT resultid="2061" eventid="19" swimtime="00:00:47.26" lane="7" heatid="19016" />
                <RESULT resultid="2060" eventid="25" swimtime="00:00:39.95" lane="4" heatid="25024" />
                <RESULT resultid="2059" eventid="37" swimtime="00:03:09.79" lane="2" heatid="37002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:34.85" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="427" birthdate="2015-01-01" gender="M" lastname="Pfeifer" firstname="Elias" license="463789">
              <RESULTS>
                <RESULT resultid="2067" eventid="20" swimtime="00:01:08.49" lane="1" heatid="20002" />
                <RESULT resultid="2066" eventid="26" swimtime="00:00:59.87" lane="4" heatid="26006" />
                <RESULT resultid="2065" eventid="30" swimtime="00:00:57.37" lane="4" heatid="30002" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="428" birthdate="2014-01-01" gender="F" lastname="Wilde" firstname="Eleonora" license="452110">
              <RESULTS>
                <RESULT resultid="2072" eventid="17" swimtime="00:01:09.40" lane="3" heatid="17009" />
                <RESULT resultid="2071" eventid="19" swimtime="00:00:59.03" lane="6" heatid="19006" />
                <RESULT resultid="2070" eventid="21" swimtime="00:01:13.65" lane="4" heatid="21006" />
                <RESULT resultid="2069" eventid="27" swimtime="00:01:05.47" lane="2" heatid="27006" />
                <RESULT resultid="2068" eventid="29" swimtime="00:00:55.37" lane="7" heatid="29004" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="429" birthdate="2015-01-01" gender="F" lastname="Rex" firstname="Caroline" license="453989">
              <RESULTS>
                <RESULT resultid="2077" eventid="17" swimtime="00:01:01.17" lane="5" heatid="17011" />
                <RESULT resultid="2076" eventid="19" swimtime="00:01:04.22" lane="3" heatid="19005" />
                <RESULT resultid="2075" eventid="25" swimtime="00:00:50.93" lane="2" heatid="25012" />
                <RESULT resultid="2074" eventid="27" swimtime="00:01:09.23" lane="2" heatid="27005" />
                <RESULT resultid="2073" eventid="29" swimtime="00:00:50.98" lane="2" heatid="29007" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="430" birthdate="2015-01-01" gender="F" lastname="Dittrich" firstname="Carolin" license="464959">
              <RESULTS>
                <RESULT resultid="2081" eventid="17" swimtime="00:01:16.15" lane="5" heatid="17002" />
                <RESULT resultid="2080" eventid="21" swimtime="00:01:23.95" lane="4" heatid="21002" />
                <RESULT resultid="2079" eventid="25" status="DNS" swimtime="00:00:00.00" lane="4" heatid="25003" />
                <RESULT resultid="2078" eventid="29" status="DNS" swimtime="00:00:00.00" lane="8" heatid="29002" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="431" birthdate="2014-01-01" gender="M" lastname="Leilich" firstname="Carl Benjamin" license="452058">
              <RESULTS>
                <RESULT resultid="2086" eventid="18" status="WDR" swimtime="00:00:00.00" lane="1" heatid="18007" />
                <RESULT resultid="2085" eventid="20" status="WDR" swimtime="00:00:00.00" lane="3" heatid="20001" />
                <RESULT resultid="2084" eventid="22" status="WDR" swimtime="00:00:00.00" lane="1" heatid="22003" />
                <RESULT resultid="2083" eventid="30" status="WDR" swimtime="00:00:00.00" lane="7" heatid="30003" />
                <RESULT resultid="2082" eventid="34" status="WDR" swimtime="00:00:00.00" lane="7" heatid="34001" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="432" birthdate="2011-01-01" gender="M" lastname="Riabtsev" firstname="Artemii" license="464433">
              <RESULTS>
                <RESULT resultid="2092" eventid="11" swimtime="00:01:33.05" lane="5" heatid="11006" />
                <RESULT resultid="2091" eventid="13" swimtime="00:00:37.26" lane="1" heatid="13006" />
                <RESULT resultid="2090" eventid="20" swimtime="00:00:51.06" lane="4" heatid="20010" />
                <RESULT resultid="2089" eventid="26" swimtime="00:00:43.21" lane="8" heatid="26018" />
                <RESULT resultid="2088" eventid="34" swimtime="00:01:23.28" lane="8" heatid="34006" />
                <RESULT resultid="2087" eventid="38" swimtime="00:03:19.21" lane="8" heatid="38002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:38.15" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="433" birthdate="2014-01-01" gender="F" lastname="Schneider" firstname="Anneta" license="459678">
              <RESULTS>
                <RESULT resultid="2097" eventid="19" swimtime="00:00:56.50" lane="5" heatid="19007" />
                <RESULT resultid="2096" eventid="21" swimtime="00:01:01.20" lane="1" heatid="21007" />
                <RESULT resultid="2095" eventid="25" swimtime="00:00:51.39" lane="1" heatid="25011" />
                <RESULT resultid="2094" eventid="29" swimtime="00:00:51.07" lane="1" heatid="29006" />
                <RESULT resultid="2093" eventid="33" swimtime="00:01:58.17" lane="1" heatid="33002" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="434" birthdate="2010-01-01" gender="F" lastname="Kunze" firstname="Anna Frida" license="426677">
              <RESULTS>
                <RESULT resultid="2101" eventid="19" swimtime="00:00:53.86" lane="8" heatid="19017" />
                <RESULT resultid="2100" eventid="23" swimtime="00:03:16.04" lane="4" heatid="23002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:34.23" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="2099" eventid="25" swimtime="00:00:44.29" lane="5" heatid="25023" />
                <RESULT resultid="2098" eventid="33" swimtime="00:01:31.52" lane="2" heatid="33009" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="435" birthdate="2010-01-01" gender="F" lastname="Bing" firstname="Adele" license="410622">
              <RESULTS>
                <RESULT resultid="2105" eventid="19" swimtime="00:00:49.70" lane="3" heatid="19017" />
                <RESULT resultid="2104" eventid="23" swimtime="00:03:16.57" lane="1" heatid="23001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:27.72" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="2103" eventid="25" swimtime="00:00:41.22" lane="4" heatid="25029" />
                <RESULT resultid="2102" eventid="33" swimtime="00:01:22.93" lane="1" heatid="33010" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
      </CLUBS>
    </MEET>
  </MEETS>
</LENEX>
