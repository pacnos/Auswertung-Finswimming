<?xml version="1.0" encoding="UTF-8"?>
<LENEX version="3.0">
  <CONSTRUCTOR name="SPLASH Meet Manager 11" registration="Nederlandse Onderwatersport Bond" version="11.77033">
    <CONTACT name="Splash Software GmbH" street="Ahornweg 41" city="Spiegel b. Bern" zip="3095" country="CH" email="sales@swimrankings.net" internet="https://www.swimrankings.net" />
  </CONSTRUCTOR>
  <MEETS>
    <MEET city="Eindhoven" name="Open NK Vinzwemmen 2023" course="LCM" deadline="2023-06-04" number="1" startmethod="1" timing="AUTOMATIC" state="NB" nation="NED">
      <AGEDATE value="2023-01-01" type="YEAR" />
      <POOL name="Pieter van den Hoogenband Zwemstadion" lanemax="9" />
      <FACILITY city="Eindhoven" name="Pieter van den Hoogenband Zwemstadion" nation="NED" state="NB" />
      <POINTTABLE pointtableid="111" name="NOB Vinzwemmen" version="2023" />
      <FEES>
        <FEE currency="EUR" type="ATHLETE" value="4500" />
      </FEES>
      <QUALIFY from="2022-01-01" until="2023-06-10" />
      <CONTACT email="nkvinzwemmen@yahoo.com" name="Karin Neehus" />
      <SESSIONS>
        <SESSION date="2023-06-24" daytime="11:45" endtime="17:00" name="Open NK Vinzwemmen ZATERDAG" number="1" officialmeeting="11:15" teamleadermeeting="10:45" warmupfrom="10:30" warmupuntil="11:15">
          <POOL lanemax="8" />
          <EVENTS>
            <EVENT eventid="1053" daytime="11:45" gender="F" number="1" order="2" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="SURFACE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1054" agemax="11" agemin="1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="29269" />
                    <RANKING order="2" place="2" resultid="28489" />
                    <RANKING order="3" place="3" resultid="29280" />
                    <RANKING order="4" place="4" resultid="28292" />
                    <RANKING order="5" place="5" resultid="28240" />
                    <RANKING order="6" place="-1" resultid="29317" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1060" agemax="13" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="28149" />
                    <RANKING order="2" place="2" resultid="29286" />
                    <RANKING order="3" place="3" resultid="28736" />
                    <RANKING order="4" place="4" resultid="29081" />
                    <RANKING order="5" place="5" resultid="28261" />
                    <RANKING order="6" place="6" resultid="28272" />
                    <RANKING order="7" place="7" resultid="28278" />
                    <RANKING order="8" place="8" resultid="29310" />
                    <RANKING order="9" place="9" resultid="29189" />
                    <RANKING order="10" place="-1" resultid="28732" />
                    <RANKING order="11" place="-1" resultid="29274" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1076" agemax="15" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="28708" />
                    <RANKING order="2" place="2" resultid="28714" />
                    <RANKING order="3" place="3" resultid="29264" />
                    <RANKING order="4" place="4" resultid="29229" />
                    <RANKING order="5" place="5" resultid="28740" />
                    <RANKING order="6" place="6" resultid="28509" />
                    <RANKING order="7" place="7" resultid="28499" />
                    <RANKING order="8" place="8" resultid="28504" />
                    <RANKING order="9" place="9" resultid="28253" />
                    <RANKING order="10" place="10" resultid="28494" />
                    <RANKING order="11" place="11" resultid="29069" />
                    <RANKING order="12" place="12" resultid="28154" />
                    <RANKING order="13" place="13" resultid="28130" />
                    <RANKING order="14" place="14" resultid="29303" />
                    <RANKING order="15" place="15" resultid="28247" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1077" agemax="17" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="28443" />
                    <RANKING order="2" place="2" resultid="29094" />
                    <RANKING order="3" place="-1" resultid="29185" />
                    <RANKING order="4" place="-1" resultid="29197" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1078" agemax="34" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="28937" />
                    <RANKING order="2" place="2" resultid="28483" />
                    <RANKING order="3" place="3" resultid="29065" />
                    <RANKING order="4" place="4" resultid="28833" />
                    <RANKING order="5" place="5" resultid="28515" />
                    <RANKING order="6" place="6" resultid="28520" />
                    <RANKING order="7" place="7" resultid="28228" />
                    <RANKING order="8" place="8" resultid="29292" />
                    <RANKING order="9" place="9" resultid="29363" />
                    <RANKING order="10" place="10" resultid="29298" />
                    <RANKING order="11" place="11" resultid="29088" />
                    <RANKING order="12" place="12" resultid="28185" />
                    <RANKING order="13" place="13" resultid="28283" />
                    <RANKING order="14" place="14" resultid="29343" />
                    <RANKING order="15" place="15" resultid="28198" />
                    <RANKING order="16" place="16" resultid="29091" />
                    <RANKING order="17" place="17" resultid="28133" />
                    <RANKING order="18" place="18" resultid="28451" />
                    <RANKING order="19" place="-1" resultid="28792" />
                    <RANKING order="20" place="-1" resultid="28106" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="12213" agemax="49" agemin="35" />
                <AGEGROUP agegroupid="1075" agemax="98" agemin="50" />
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="1079" daytime="12:00" gender="M" number="2" order="3" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="SURFACE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1080" agemax="11" agemin="1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="29100" />
                    <RANKING order="2" place="2" resultid="28159" />
                    <RANKING order="3" place="3" resultid="29360" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1081" agemax="13" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="28525" />
                    <RANKING order="2" place="2" resultid="29336" />
                    <RANKING order="3" place="3" resultid="28761" />
                    <RANKING order="4" place="4" resultid="29117" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1082" agemax="15" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="29224" />
                    <RANKING order="2" place="2" resultid="29110" />
                    <RANKING order="3" place="3" resultid="28728" />
                    <RANKING order="4" place="4" resultid="29239" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1083" agemax="17" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="28691" />
                    <RANKING order="2" place="2" resultid="28852" />
                    <RANKING order="3" place="3" resultid="28530" />
                    <RANKING order="4" place="4" resultid="29104" />
                    <RANKING order="5" place="5" resultid="28212" />
                    <RANKING order="6" place="-1" resultid="29201" />
                    <RANKING order="7" place="-1" resultid="29193" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1084" agemax="34" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="28787" />
                    <RANKING order="2" place="2" resultid="28796" />
                    <RANKING order="3" place="3" resultid="28724" />
                    <RANKING order="4" place="4" resultid="28686" />
                    <RANKING order="5" place="5" resultid="29205" />
                    <RANKING order="6" place="6" resultid="28172" />
                    <RANKING order="7" place="7" resultid="29214" />
                    <RANKING order="8" place="8" resultid="28535" />
                    <RANKING order="9" place="9" resultid="29216" />
                    <RANKING order="10" place="10" resultid="28232" />
                    <RANKING order="11" place="11" resultid="28843" />
                    <RANKING order="12" place="12" resultid="28460" />
                    <RANKING order="13" place="13" resultid="28179" />
                    <RANKING order="14" place="14" resultid="28164" />
                    <RANKING order="15" place="15" resultid="28117" />
                    <RANKING order="16" place="16" resultid="29369" />
                    <RANKING order="17" place="-1" resultid="28473" />
                    <RANKING order="18" place="-1" resultid="28191" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="12214" agemax="49" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="28846" />
                    <RANKING order="2" place="2" resultid="28219" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1085" agemax="98" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="29351" />
                    <RANKING order="2" place="2" resultid="28205" />
                    <RANKING order="3" place="3" resultid="29329" />
                    <RANKING order="4" place="4" resultid="28111" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="1093" daytime="12:15" gender="F" number="3" order="4" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="1500" relaycount="1" stroke="SURFACE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1095" agemax="13" agemin="12" />
                <AGEGROUP agegroupid="29415" agemax="15" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="28703" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1096" agemax="17" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="29219" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="29417" agemax="34" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="29260" />
                    <RANKING order="2" place="2" resultid="28452" />
                    <RANKING order="3" place="3" resultid="29092" />
                    <RANKING order="4" place="4" resultid="28142" />
                    <RANKING order="5" place="5" resultid="29089" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="12215" agemax="49" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="28268" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1098" agemax="98" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="28435" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="18215" daytime="13:00" gender="M" number="4" order="6" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="1500" relaycount="1" stroke="SURFACE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="18216" agemax="13" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="29467" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="18217" agemax="15" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="29463" />
                    <RANKING order="2" place="2" resultid="29468" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="18218" agemax="17" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="29465" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="18219" agemax="34" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="29464" />
                    <RANKING order="2" place="2" resultid="29462" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="18220" agemax="49" agemin="35" />
                <AGEGROUP agegroupid="18221" agemax="98" agemin="50" />
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="22849" daytime="13:25" gender="F" number="5" order="7" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="800" relaycount="1" stroke="IMMERSION" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="22851" agemax="15" agemin="14" />
                <AGEGROUP agegroupid="22852" agemax="17" agemin="16" />
                <AGEGROUP agegroupid="22853" agemax="34" agemin="18" />
                <AGEGROUP agegroupid="22854" agemax="49" agemin="35" />
                <AGEGROUP agegroupid="22855" agemax="98" agemin="50" />
                <AGEGROUP agegroupid="23121" agemax="15" agemin="14" />
                <AGEGROUP agegroupid="23134" agemax="17" agemin="16" />
                <AGEGROUP agegroupid="24839" agemax="34" agemin="18" />
                <AGEGROUP agegroupid="24840" agemax="49" agemin="35" />
                <AGEGROUP agegroupid="23136" agemax="98" agemin="50" />
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="26746" daytime="13:25" number="6" order="9" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="800" relaycount="1" stroke="IMMERSION" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="26747" agemax="15" agemin="14" gender="M" />
                <AGEGROUP agegroupid="26748" agemax="17" agemin="16" gender="M">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="29249" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="26749" agemax="34" agemin="18" gender="M">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="28173" />
                    <RANKING order="2" place="2" resultid="29255" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="26750" agemax="49" agemin="35" gender="M" />
                <AGEGROUP agegroupid="26751" agemax="98" agemin="50" gender="M" />
                <AGEGROUP agegroupid="29433" agemax="34" agemin="18" gender="F">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="29434" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="7254" daytime="13:35" gender="F" number="7" order="10" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BIFINS" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="8048" agemax="11" agemin="1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="28293" />
                    <RANKING order="2" place="2" resultid="29318" />
                    <RANKING order="3" place="3" resultid="28241" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7255" agemax="13" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="28273" />
                    <RANKING order="2" place="2" resultid="28262" />
                    <RANKING order="3" place="3" resultid="29311" />
                    <RANKING order="4" place="-1" resultid="29190" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7256" agemax="15" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="29230" />
                    <RANKING order="2" place="2" resultid="29070" />
                    <RANKING order="3" place="3" resultid="28254" />
                    <RANKING order="4" place="4" resultid="28155" />
                    <RANKING order="5" place="5" resultid="29304" />
                    <RANKING order="6" place="6" resultid="28248" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7257" agemax="17" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="29164" />
                    <RANKING order="2" place="2" resultid="28444" />
                    <RANKING order="3" place="3" resultid="29442" />
                    <RANKING order="4" place="4" resultid="29186" />
                    <RANKING order="5" place="5" resultid="29198" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7258" agemax="34" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="29150" />
                    <RANKING order="2" place="2" resultid="29446" />
                    <RANKING order="3" place="3" resultid="28186" />
                    <RANKING order="4" place="4" resultid="28284" />
                    <RANKING order="5" place="5" resultid="28199" />
                    <RANKING order="6" place="6" resultid="29344" />
                    <RANKING order="7" place="7" resultid="28134" />
                    <RANKING order="8" place="8" resultid="28143" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="12218" agemax="49" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="28269" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7259" agemax="98" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="28436" />
                    <RANKING order="2" place="2" resultid="29158" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="7271" daytime="13:55" gender="M" number="8" order="11" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BIFINS" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="8049" agemax="11" agemin="1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="28160" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7272" agemax="13" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="29337" />
                    <RANKING order="2" place="2" resultid="28762" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7273" agemax="15" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="29154" />
                    <RANKING order="2" place="2" resultid="29077" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7274" agemax="17" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="28836" />
                    <RANKING order="2" place="2" resultid="28213" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7275" agemax="34" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="28800" />
                    <RANKING order="2" place="2" resultid="29217" />
                    <RANKING order="3" place="3" resultid="28118" />
                    <RANKING order="4" place="4" resultid="28192" />
                    <RANKING order="5" place="5" resultid="29172" />
                    <RANKING order="6" place="6" resultid="28180" />
                    <RANKING order="7" place="7" resultid="28165" />
                    <RANKING order="8" place="8" resultid="28461" />
                    <RANKING order="9" place="9" resultid="29162" />
                    <RANKING order="10" place="10" resultid="29370" />
                    <RANKING order="11" place="-1" resultid="28101" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="12219" agemax="49" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="28220" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7276" agemax="98" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="29352" />
                    <RANKING order="2" place="2" resultid="28206" />
                    <RANKING order="3" place="3" resultid="28112" />
                    <RANKING order="4" place="4" resultid="29330" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="26758" daytime="14:10" gender="F" number="9" order="13" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="SURFACE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="26759" agemax="11" agemin="1" calculate="TOTAL" />
                <AGEGROUP agegroupid="26760" agemax="13" agemin="12" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="28298" />
                    <RANKING order="2" place="2" resultid="29381" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="26761" agemax="15" agemin="14" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="29388" />
                    <RANKING order="2" place="2" resultid="29486" />
                    <RANKING order="3" place="3" resultid="28540" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="26762" agemax="17" agemin="16" calculate="TOTAL" />
                <AGEGROUP agegroupid="26763" agemax="34" agemin="18" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="29379" />
                    <RANKING order="2" place="2" resultid="29386" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="26764" agemax="49" agemin="35" calculate="TOTAL" />
                <AGEGROUP agegroupid="26765" agemax="98" agemin="50" calculate="TOTAL" />
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="26768" daytime="14:20" gender="M" number="10" order="14" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="SURFACE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="26769" agemax="11" agemin="1" calculate="TOTAL" />
                <AGEGROUP agegroupid="26770" agemax="13" agemin="12" calculate="TOTAL" />
                <AGEGROUP agegroupid="26771" agemax="15" agemin="14" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="29390" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="26772" agemax="17" agemin="16" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="29122" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="26773" agemax="34" agemin="18" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="29244" />
                    <RANKING order="2" place="2" resultid="29473" />
                    <RANKING order="3" place="3" resultid="29481" />
                    <RANKING order="4" place="-1" resultid="29389" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="26774" agemax="49" agemin="35" calculate="TOTAL" />
                <AGEGROUP agegroupid="26775" agemax="98" agemin="50" calculate="TOTAL" />
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="1120" daytime="15:10" gender="F" number="11" order="16" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BIFINS" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1121" agemax="11" agemin="1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="29319" />
                    <RANKING order="2" place="2" resultid="28294" />
                    <RANKING order="3" place="3" resultid="28242" />
                    <RANKING order="4" place="3" resultid="29281" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1122" agemax="13" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="29074" />
                    <RANKING order="2" place="2" resultid="28263" />
                    <RANKING order="3" place="3" resultid="28274" />
                    <RANKING order="4" place="4" resultid="29275" />
                    <RANKING order="5" place="5" resultid="29312" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1123" agemax="15" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="28741" />
                    <RANKING order="2" place="2" resultid="28156" />
                    <RANKING order="3" place="3" resultid="28255" />
                    <RANKING order="4" place="4" resultid="29305" />
                    <RANKING order="5" place="5" resultid="28131" />
                    <RANKING order="6" place="6" resultid="28249" />
                    <RANKING order="7" place="-1" resultid="29231" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1124" agemax="17" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="29165" />
                    <RANKING order="2" place="-1" resultid="29441" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1125" agemax="34" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="28938" />
                    <RANKING order="2" place="2" resultid="29151" />
                    <RANKING order="3" place="3" resultid="28793" />
                    <RANKING order="4" place="4" resultid="29066" />
                    <RANKING order="5" place="5" resultid="29445" />
                    <RANKING order="6" place="6" resultid="29364" />
                    <RANKING order="7" place="7" resultid="28187" />
                    <RANKING order="8" place="8" resultid="28135" />
                    <RANKING order="9" place="9" resultid="28200" />
                    <RANKING order="10" place="10" resultid="28144" />
                    <RANKING order="11" place="11" resultid="28285" />
                    <RANKING order="12" place="12" resultid="28453" />
                    <RANKING order="13" place="13" resultid="28107" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="12220" agemax="49" agemin="35" />
                <AGEGROUP agegroupid="1126" agemax="98" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="29159" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="1127" daytime="15:15" gender="M" number="12" order="17" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BIFINS" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1128" agemax="11" agemin="1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="28161" />
                    <RANKING order="2" place="2" resultid="29361" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1129" agemax="13" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="29338" />
                    <RANKING order="2" place="2" resultid="28767" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1130" agemax="15" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="29155" />
                    <RANKING order="2" place="2" resultid="29225" />
                    <RANKING order="3" place="3" resultid="29079" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1131" agemax="17" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="28837" />
                    <RANKING order="2" place="2" resultid="29194" />
                    <RANKING order="3" place="3" resultid="28214" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1132" agemax="34" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="28801" />
                    <RANKING order="2" place="2" resultid="29443" />
                    <RANKING order="3" place="3" resultid="28844" />
                    <RANKING order="4" place="4" resultid="29215" />
                    <RANKING order="5" place="5" resultid="28102" />
                    <RANKING order="6" place="6" resultid="29206" />
                    <RANKING order="7" place="7" resultid="29218" />
                    <RANKING order="8" place="8" resultid="28840" />
                    <RANKING order="9" place="9" resultid="28234" />
                    <RANKING order="10" place="10" resultid="28119" />
                    <RANKING order="11" place="11" resultid="28462" />
                    <RANKING order="12" place="12" resultid="28181" />
                    <RANKING order="13" place="13" resultid="29173" />
                    <RANKING order="14" place="14" resultid="28193" />
                    <RANKING order="15" place="15" resultid="29371" />
                    <RANKING order="16" place="16" resultid="29163" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="12221" agemax="49" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="28221" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1133" agemax="98" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="29353" />
                    <RANKING order="2" place="2" resultid="28207" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="7278" daytime="15:25" gender="F" number="13" order="18" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="SURFACE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="8050" agemax="11" agemin="1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="29270" />
                    <RANKING order="2" place="2" resultid="28490" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7279" agemax="13" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="28150" />
                    <RANKING order="2" place="2" resultid="28737" />
                    <RANKING order="3" place="3" resultid="29287" />
                    <RANKING order="4" place="4" resultid="28733" />
                    <RANKING order="5" place="5" resultid="28279" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7280" agemax="15" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="28715" />
                    <RANKING order="2" place="2" resultid="28704" />
                    <RANKING order="3" place="3" resultid="28500" />
                    <RANKING order="4" place="4" resultid="29235" />
                    <RANKING order="5" place="5" resultid="28510" />
                    <RANKING order="6" place="6" resultid="28505" />
                    <RANKING order="7" place="7" resultid="28495" />
                    <RANKING order="8" place="8" resultid="28157" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7281" agemax="17" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="29220" />
                    <RANKING order="2" place="2" resultid="28445" />
                    <RANKING order="3" place="3" resultid="29095" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7282" agemax="34" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="28479" />
                    <RANKING order="2" place="2" resultid="28484" />
                    <RANKING order="3" place="3" resultid="28516" />
                    <RANKING order="4" place="4" resultid="28521" />
                    <RANKING order="5" place="5" resultid="29090" />
                    <RANKING order="6" place="6" resultid="28454" />
                    <RANKING order="7" place="7" resultid="29299" />
                    <RANKING order="8" place="8" resultid="29293" />
                    <RANKING order="9" place="9" resultid="29093" />
                    <RANKING order="10" place="10" resultid="28286" />
                    <RANKING order="11" place="11" resultid="29345" />
                    <RANKING order="12" place="12" resultid="28136" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="12222" agemax="49" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="28270" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7283" agemax="98" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="28437" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="7264" daytime="15:50" gender="M" number="14" order="20" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="SURFACE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="7265" agemax="11" agemin="1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="28162" />
                    <RANKING order="2" place="2" resultid="29101" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8643" agemax="13" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="28526" />
                    <RANKING order="2" place="2" resultid="29119" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7266" agemax="15" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="28698" />
                    <RANKING order="2" place="2" resultid="28729" />
                    <RANKING order="3" place="3" resultid="29112" />
                    <RANKING order="4" place="-1" resultid="29240" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7267" agemax="17" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="28853" />
                    <RANKING order="2" place="2" resultid="29250" />
                    <RANKING order="3" place="3" resultid="28531" />
                    <RANKING order="4" place="4" resultid="29105" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7268" agemax="34" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="28788" />
                    <RANKING order="2" place="2" resultid="28687" />
                    <RANKING order="3" place="3" resultid="28235" />
                    <RANKING order="4" place="4" resultid="28166" />
                    <RANKING order="5" place="5" resultid="28120" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="12223" agemax="49" agemin="35" />
                <AGEGROUP agegroupid="7269" agemax="98" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="29331" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="1105" daytime="16:10" gender="F" number="15" order="21" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="IMMERSION" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1106" agemax="13" agemin="12" />
                <AGEGROUP agegroupid="1107" agemax="15" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="29265" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1108" agemax="17" agemin="16" />
                <AGEGROUP agegroupid="1109" agemax="34" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="28145" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="12224" agemax="49" agemin="35" />
                <AGEGROUP agegroupid="1110" agemax="98" agemin="50" />
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="1114" daytime="16:20" gender="M" number="16" order="22" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="IMMERSION" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1115" agemax="13" agemin="12" />
                <AGEGROUP agegroupid="1116" agemax="15" agemin="14" />
                <AGEGROUP agegroupid="1117" agemax="17" agemin="16" />
                <AGEGROUP agegroupid="1118" agemax="34" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="28474" />
                    <RANKING order="2" place="2" resultid="29256" />
                    <RANKING order="3" place="3" resultid="28725" />
                    <RANKING order="4" place="4" resultid="28174" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="12225" agemax="49" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="28847" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1119" agemax="98" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="28113" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="1140" daytime="16:40" gender="X" number="17" order="25" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="4" stroke="BIFINS" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="28544" agemax="11" agemin="1" calculate="TOTAL" />
                <AGEGROUP agegroupid="28545" agemax="13" agemin="12" />
                <AGEGROUP agegroupid="28546" agemax="15" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="29391" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="28547" agemax="17" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="29392" />
                    <RANKING order="2" place="2" resultid="29210" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="28548" agemax="34" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="29489" />
                    <RANKING order="2" place="2" resultid="29176" />
                    <RANKING order="3" place="3" resultid="29482" />
                    <RANKING order="4" place="4" resultid="29490" />
                    <RANKING order="5" place="5" resultid="28177" />
                    <RANKING order="6" place="6" resultid="29384" />
                    <RANKING order="7" place="7" resultid="29488" />
                    <RANKING order="8" place="-1" resultid="29245" />
                    <RANKING order="9" place="-1" resultid="29385" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="28549" agemax="49" agemin="35" />
                <AGEGROUP agegroupid="28550" agemax="98" agemin="50" />
              </AGEGROUPS>
            </EVENT>
          </EVENTS>
          <JUDGES>
            <JUDGE officialid="2149" remarks="ok" />
            <JUDGE officialid="21300" remarks="ok" />
            <JUDGE officialid="21329" remarks="ok" />
            <JUDGE officialid="24070" remarks="ok" />
            <JUDGE officialid="28781" remarks="ok" />
            <JUDGE officialid="1520" remarks="ok" />
            <JUDGE officialid="25526" remarks="ok" />
            <JUDGE officialid="1510" remarks="ok" />
            <JUDGE officialid="6661" remarks="ok" />
            <JUDGE officialid="28777" remarks="ok" />
            <JUDGE officialid="7858" remarks="ok" />
            <JUDGE officialid="21127" remarks="ok" />
            <JUDGE officialid="2140" remarks="ok" />
            <JUDGE officialid="21335" remarks="ok" />
            <JUDGE officialid="26602" remarks="ok" />
            <JUDGE officialid="1538" remarks="ok" />
            <JUDGE officialid="29057" remarks="ok" />
            <JUDGE number="101" officialid="4863" remarks="ok" />
            <JUDGE number="102" officialid="28783" remarks="ok" />
            <JUDGE number="103" officialid="2781" remarks="ok" />
            <JUDGE number="104" officialid="23071" remarks="ok" />
            <JUDGE number="204" officialid="28487" remarks="ok" />
            <JUDGE number="105" officialid="2148" remarks="ok" />
            <JUDGE number="106" officialid="5128" remarks="ok" />
            <JUDGE number="107" officialid="25528" remarks="ok" />
            <JUDGE number="108" officialid="27674" remarks="ok" />
            <JUDGE officialid="25527" remarks="reserve" />
            <JUDGE number="1" officialid="6383" remarks="OCEANUS" />
            <JUDGE number="2" officialid="3072" remarks="Orka &apos;97" />
            <JUDGE number="3" officialid="4401" remarks="OSV Delphis en Emese" />
            <JUDGE number="4" officialid="3074" remarks="OWT PONTOS en Mahmoud" />
            <JUDGE number="5" officialid="3073" remarks="VZ Utrecht" />
            <JUDGE number="6" officialid="27676" remarks="Waves" />
            <JUDGE number="7" officialid="1536" remarks="MonoVinzz" />
            <JUDGE number="8" officialid="24198" remarks="DJK-VfR Muhlheim" />
            <JUDGE number="9" officialid="24196" remarks="TC Heilbronn" />
            <JUDGE number="10" officialid="24200" remarks="CS Gravenchon" />
            <JUDGE number="11" officialid="28804" remarks="SC DHfK Leipzig" />
            <JUDGE number="12" officialid="28804" remarks="TC Delitzsch" />
            <JUDGE number="13" officialid="28803" remarks="1. Chemnitz TVeV" />
            <JUDGE number="14" officialid="29436" remarks="Swiss Team" />
            <JUDGE number="15" officialid="27686" remarks="TC Nemo Plauen" />
            <JUDGE number="16" officialid="27807" remarks="PF NAP Aix" />
            <JUDGE number="17" officialid="28824" remarks="CSA Kremlin Bicetre" />
            <JUDGE number="18" officialid="24572" remarks="Tours NAP" />
            <JUDGE number="19" officialid="24482" remarks="Club Ciotaden NP" />
            <JUDGE number="20" officialid="27826" remarks="CPB NAP" />
            <JUDGE number="21" officialid="27683" remarks="Binger TSCeV" />
            <JUDGE number="22" officialid="24196" remarks="TC Harz" />
            <JUDGE number="23" officialid="24569" remarks="TC fez Berlin" />
            <JUDGE number="24" officialid="29179" remarks="LGM" />
            <JUDGE number="25" officialid="24573" remarks="Nautilus" />
            <JUDGE number="26" officialid="24795" remarks="Aq-Nivelles" />
          </JUDGES>
        </SESSION>
        <SESSION date="2023-06-25" daytime="11:15" endtime="16:12" name="Open NK Vinzwemmen ZONDAG" number="2" officialmeeting="10:45" teamleadermeeting="10:30" warmupfrom="10:30" warmupuntil="11:15">
          <POOL lanemin="1" lanemax="8" />
          <EVENTS>
            <EVENT eventid="1147" daytime="11:15" gender="F" number="18" order="2" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="APNEA" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1149" agemax="15" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="28709" />
                    <RANKING order="2" place="2" resultid="29266" />
                    <RANKING order="3" place="3" resultid="29232" />
                    <RANKING order="4" place="4" resultid="28511" />
                    <RANKING order="5" place="5" resultid="28742" />
                    <RANKING order="6" place="6" resultid="28501" />
                    <RANKING order="7" place="7" resultid="28506" />
                    <RANKING order="8" place="8" resultid="28256" />
                    <RANKING order="9" place="9" resultid="28496" />
                    <RANKING order="10" place="10" resultid="28468" />
                    <RANKING order="11" place="11" resultid="29071" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1150" agemax="17" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="28446" />
                    <RANKING order="2" place="2" resultid="29096" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1151" agemax="34" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="28939" />
                    <RANKING order="2" place="2" resultid="28794" />
                    <RANKING order="3" place="3" resultid="28480" />
                    <RANKING order="4" place="4" resultid="28485" />
                    <RANKING order="5" place="5" resultid="28834" />
                    <RANKING order="6" place="6" resultid="29067" />
                    <RANKING order="7" place="7" resultid="28517" />
                    <RANKING order="8" place="8" resultid="28522" />
                    <RANKING order="9" place="9" resultid="28229" />
                    <RANKING order="10" place="10" resultid="29300" />
                    <RANKING order="11" place="11" resultid="28287" />
                    <RANKING order="12" place="12" resultid="29346" />
                    <RANKING order="13" place="13" resultid="29365" />
                    <RANKING order="14" place="14" resultid="28126" />
                    <RANKING order="15" place="15" resultid="28108" />
                    <RANKING order="16" place="16" resultid="28201" />
                    <RANKING order="17" place="-1" resultid="28455" />
                    <RANKING order="18" place="-1" resultid="29294" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="12228" agemax="49" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="29324" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1152" agemax="98" agemin="50" />
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="1153" daytime="11:25" gender="M" number="19" order="3" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="APNEA" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1154" agemax="15" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="29226" />
                    <RANKING order="2" place="-1" resultid="29241" />
                    <RANKING order="3" place="-1" resultid="29113" />
                    <RANKING order="4" place="-1" resultid="29156" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1155" agemax="17" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="28532" />
                    <RANKING order="2" place="2" resultid="28693" />
                    <RANKING order="3" place="3" resultid="29106" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1156" agemax="34" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="28475" />
                    <RANKING order="2" place="2" resultid="28789" />
                    <RANKING order="3" place="3" resultid="28536" />
                    <RANKING order="4" place="4" resultid="29207" />
                    <RANKING order="5" place="5" resultid="28688" />
                    <RANKING order="6" place="6" resultid="28463" />
                    <RANKING order="7" place="7" resultid="28845" />
                    <RANKING order="8" place="8" resultid="28236" />
                    <RANKING order="9" place="9" resultid="28121" />
                    <RANKING order="10" place="10" resultid="28194" />
                    <RANKING order="11" place="11" resultid="28167" />
                    <RANKING order="12" place="12" resultid="29372" />
                    <RANKING order="13" place="-1" resultid="28797" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="12229" agemax="49" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="28848" />
                    <RANKING order="2" place="2" resultid="28222" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1157" agemax="98" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="29354" />
                    <RANKING order="2" place="2" resultid="29332" />
                    <RANKING order="3" place="3" resultid="28208" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="1158" daytime="11:35" gender="F" number="20" order="4" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="800" relaycount="1" stroke="SURFACE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="26270" agemax="13" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="28738" />
                    <RANKING order="2" place="2" resultid="28734" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="16171" agemax="15" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="28705" />
                    <RANKING order="2" place="2" resultid="29233" />
                    <RANKING order="3" place="3" resultid="28512" />
                    <RANKING order="4" place="4" resultid="29236" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="16172" agemax="17" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="29221" />
                    <RANKING order="2" place="2" resultid="29097" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="16173" agemax="34" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="29261" />
                    <RANKING order="2" place="2" resultid="28456" />
                    <RANKING order="3" place="3" resultid="28288" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="16174" agemax="49" agemin="35" />
                <AGEGROUP agegroupid="16175" agemax="98" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="28438" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="16574" daytime="12:00" gender="M" number="21" order="5" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="800" relaycount="1" stroke="SURFACE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="26020" agemax="13" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="28527" />
                    <RANKING order="2" place="2" resultid="29120" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="16575" agemax="15" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="28699" />
                    <RANKING order="2" place="2" resultid="28730" />
                    <RANKING order="3" place="3" resultid="29114" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="16577" agemax="17" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="28854" />
                    <RANKING order="2" place="2" resultid="29251" />
                    <RANKING order="3" place="3" resultid="29107" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="16579" agemax="34" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="28726" />
                    <RANKING order="2" place="2" resultid="28175" />
                    <RANKING order="3" place="3" resultid="29257" />
                    <RANKING order="4" place="4" resultid="29170" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="16581" agemax="49" agemin="35" />
                <AGEGROUP agegroupid="16583" agemax="98" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="28114" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="1168" daytime="12:25" gender="F" number="22" order="6" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BIFINS" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1169" agemax="11" agemin="1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="28491" />
                    <RANKING order="2" place="2" resultid="29320" />
                    <RANKING order="3" place="3" resultid="28295" />
                    <RANKING order="4" place="4" resultid="29282" />
                    <RANKING order="5" place="5" resultid="28243" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1170" agemax="13" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="29288" />
                    <RANKING order="2" place="2" resultid="29075" />
                    <RANKING order="3" place="3" resultid="28275" />
                    <RANKING order="4" place="4" resultid="28264" />
                    <RANKING order="5" place="5" resultid="28280" />
                    <RANKING order="6" place="6" resultid="29276" />
                    <RANKING order="7" place="7" resultid="29191" />
                    <RANKING order="8" place="8" resultid="29313" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1171" agemax="15" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="28469" />
                    <RANKING order="2" place="2" resultid="28257" />
                    <RANKING order="3" place="3" resultid="29306" />
                    <RANKING order="4" place="4" resultid="28250" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1172" agemax="17" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="29166" />
                    <RANKING order="2" place="2" resultid="28447" />
                    <RANKING order="3" place="3" resultid="29199" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1173" agemax="34" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="29152" />
                    <RANKING order="2" place="2" resultid="29366" />
                    <RANKING order="3" place="3" resultid="28188" />
                    <RANKING order="4" place="4" resultid="28458" />
                    <RANKING order="5" place="5" resultid="28127" />
                    <RANKING order="6" place="6" resultid="28202" />
                    <RANKING order="7" place="7" resultid="28137" />
                    <RANKING order="8" place="8" resultid="29347" />
                    <RANKING order="9" place="9" resultid="28146" />
                    <RANKING order="10" place="10" resultid="28109" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="12232" agemax="49" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="29325" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1174" agemax="98" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="28439" />
                    <RANKING order="2" place="2" resultid="29160" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="1175" daytime="12:40" gender="M" number="23" order="7" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BIFINS" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1176" agemax="11" agemin="1" />
                <AGEGROUP agegroupid="1177" agemax="13" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="29339" />
                    <RANKING order="2" place="2" resultid="28763" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1178" agemax="15" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="29078" />
                    <RANKING order="2" place="-1" resultid="29157" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1179" agemax="17" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="28838" />
                    <RANKING order="2" place="2" resultid="29202" />
                    <RANKING order="3" place="3" resultid="28215" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1180" agemax="34" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="28802" />
                    <RANKING order="2" place="2" resultid="29444" />
                    <RANKING order="3" place="3" resultid="28103" />
                    <RANKING order="4" place="4" resultid="28237" />
                    <RANKING order="5" place="5" resultid="28122" />
                    <RANKING order="6" place="6" resultid="28464" />
                    <RANKING order="7" place="7" resultid="28841" />
                    <RANKING order="8" place="8" resultid="29174" />
                    <RANKING order="9" place="9" resultid="28168" />
                    <RANKING order="10" place="10" resultid="29373" />
                    <RANKING order="11" place="11" resultid="29167" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="12233" agemax="49" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="28223" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1181" agemax="98" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="29355" />
                    <RANKING order="2" place="2" resultid="28209" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="1210" daytime="12:50" gender="X" number="24" order="9" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="APNEA" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1213" agemax="15" agemin="14" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="29246" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="26610" agemax="17" agemin="16" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="29394" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1215" agemax="34" agemin="18" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="29393" />
                    <RANKING order="2" place="2" resultid="28539" />
                    <RANKING order="3" place="3" resultid="29382" />
                    <RANKING order="4" place="4" resultid="29483" />
                    <RANKING order="5" place="5" resultid="29492" />
                    <RANKING order="6" place="6" resultid="29177" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="12240" agemax="49" agemin="35" calculate="TOTAL" />
                <AGEGROUP agegroupid="1216" agemax="98" agemin="50" calculate="TOTAL" />
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="7287" daytime="13:40" gender="F" number="25" order="11" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="SURFACE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="7288" agemax="11" agemin="1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="29271" />
                    <RANKING order="2" place="2" resultid="28492" />
                    <RANKING order="3" place="3" resultid="29283" />
                    <RANKING order="4" place="4" resultid="28296" />
                    <RANKING order="5" place="5" resultid="29321" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7289" agemax="13" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="29289" />
                    <RANKING order="2" place="2" resultid="28739" />
                    <RANKING order="3" place="3" resultid="29076" />
                    <RANKING order="4" place="4" resultid="28735" />
                    <RANKING order="5" place="5" resultid="28265" />
                    <RANKING order="6" place="6" resultid="29277" />
                    <RANKING order="7" place="7" resultid="29314" />
                    <RANKING order="8" place="8" resultid="29192" />
                    <RANKING order="9" place="-1" resultid="28151" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7290" agemax="15" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="28710" />
                    <RANKING order="2" place="2" resultid="28716" />
                    <RANKING order="3" place="3" resultid="29234" />
                    <RANKING order="4" place="4" resultid="28743" />
                    <RANKING order="5" place="5" resultid="28502" />
                    <RANKING order="6" place="6" resultid="28769" />
                    <RANKING order="7" place="7" resultid="29237" />
                    <RANKING order="8" place="8" resultid="28507" />
                    <RANKING order="9" place="9" resultid="28258" />
                    <RANKING order="10" place="10" resultid="28497" />
                    <RANKING order="11" place="11" resultid="28470" />
                    <RANKING order="12" place="12" resultid="29307" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7291" agemax="17" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="28448" />
                    <RANKING order="2" place="2" resultid="29187" />
                    <RANKING order="3" place="3" resultid="29200" />
                    <RANKING order="4" place="4" resultid="29098" />
                    <RANKING order="5" place="-1" resultid="29222" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7292" agemax="34" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="28940" />
                    <RANKING order="2" place="2" resultid="28481" />
                    <RANKING order="3" place="3" resultid="28486" />
                    <RANKING order="4" place="4" resultid="29068" />
                    <RANKING order="5" place="5" resultid="28523" />
                    <RANKING order="6" place="6" resultid="28518" />
                    <RANKING order="7" place="7" resultid="29301" />
                    <RANKING order="8" place="8" resultid="29367" />
                    <RANKING order="9" place="9" resultid="29348" />
                    <RANKING order="10" place="10" resultid="28289" />
                    <RANKING order="11" place="11" resultid="28203" />
                    <RANKING order="12" place="12" resultid="28457" />
                    <RANKING order="13" place="13" resultid="28128" />
                    <RANKING order="14" place="14" resultid="28138" />
                    <RANKING order="15" place="-1" resultid="28795" />
                    <RANKING order="16" place="-1" resultid="29295" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="12234" agemax="49" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="29326" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7293" agemax="98" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="28440" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="7295" daytime="14:00" gender="M" number="26" order="12" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="SURFACE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="7296" agemax="11" agemin="1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="29102" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7297" agemax="13" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="28528" />
                    <RANKING order="2" place="2" resultid="28764" />
                    <RANKING order="3" place="3" resultid="29340" />
                    <RANKING order="4" place="4" resultid="29121" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7298" agemax="15" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="28700" />
                    <RANKING order="2" place="2" resultid="29227" />
                    <RANKING order="3" place="3" resultid="29115" />
                    <RANKING order="4" place="4" resultid="28731" />
                    <RANKING order="5" place="-1" resultid="29242" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7299" agemax="17" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="28694" />
                    <RANKING order="2" place="2" resultid="28533" />
                    <RANKING order="3" place="3" resultid="29108" />
                    <RANKING order="4" place="4" resultid="29195" />
                    <RANKING order="5" place="5" resultid="28216" />
                    <RANKING order="6" place="-1" resultid="29203" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7300" agemax="34" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="28790" />
                    <RANKING order="2" place="2" resultid="29208" />
                    <RANKING order="3" place="3" resultid="28537" />
                    <RANKING order="4" place="4" resultid="28465" />
                    <RANKING order="5" place="5" resultid="28182" />
                    <RANKING order="6" place="6" resultid="28169" />
                    <RANKING order="7" place="7" resultid="28195" />
                    <RANKING order="8" place="8" resultid="29375" />
                    <RANKING order="9" place="-1" resultid="28476" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="12235" agemax="49" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="28224" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7301" agemax="98" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="29356" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="1196" daytime="14:15" gender="F" number="27" order="13" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="BIFINS" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1197" agemax="11" agemin="1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="28244" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1198" agemax="13" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="28276" />
                    <RANKING order="2" place="2" resultid="28281" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1199" agemax="15" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="29072" />
                    <RANKING order="2" place="2" resultid="28251" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1200" agemax="17" agemin="16" />
                <AGEGROUP agegroupid="1201" agemax="34" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="29153" />
                    <RANKING order="2" place="2" resultid="28189" />
                    <RANKING order="3" place="3" resultid="28147" />
                    <RANKING order="4" place="4" resultid="28139" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="12236" agemax="49" agemin="35" />
                <AGEGROUP agegroupid="1202" agemax="98" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="29161" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="1203" daytime="14:30" gender="M" number="28" order="14" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="BIFINS" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1204" agemax="11" agemin="1" />
                <AGEGROUP agegroupid="1205" agemax="13" agemin="12" />
                <AGEGROUP agegroupid="1206" agemax="15" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="29080" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1207" agemax="17" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="28839" />
                    <RANKING order="2" place="2" resultid="29252" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1208" agemax="34" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="28238" />
                    <RANKING order="2" place="2" resultid="28104" />
                    <RANKING order="3" place="3" resultid="29175" />
                    <RANKING order="4" place="4" resultid="29171" />
                    <RANKING order="5" place="5" resultid="28123" />
                    <RANKING order="6" place="6" resultid="29168" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="12237" agemax="49" agemin="35" />
                <AGEGROUP agegroupid="1209" agemax="98" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="28210" />
                    <RANKING order="2" place="2" resultid="29333" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="1182" daytime="14:40" gender="F" number="29" order="16" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="IMMERSION" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1183" agemax="13" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="28152" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1184" agemax="15" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="28711" />
                    <RANKING order="2" place="2" resultid="29267" />
                    <RANKING order="3" place="3" resultid="28706" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1185" agemax="17" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="28449" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1186" agemax="34" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="29485" />
                    <RANKING order="2" place="2" resultid="28835" />
                    <RANKING order="3" place="3" resultid="28519" />
                    <RANKING order="4" place="4" resultid="28524" />
                    <RANKING order="5" place="5" resultid="28230" />
                    <RANKING order="6" place="6" resultid="29349" />
                    <RANKING order="7" place="7" resultid="28148" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="12238" agemax="49" agemin="35" />
                <AGEGROUP agegroupid="1187" agemax="98" agemin="50" />
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="1190" daytime="14:50" gender="M" number="30" order="17" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="IMMERSION" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1191" agemax="13" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="28765" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1192" agemax="15" agemin="14" />
                <AGEGROUP agegroupid="1193" agemax="17" agemin="16" />
                <AGEGROUP agegroupid="1194" agemax="34" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="28791" />
                    <RANKING order="2" place="2" resultid="28798" />
                    <RANKING order="3" place="3" resultid="28727" />
                    <RANKING order="4" place="4" resultid="28538" />
                    <RANKING order="5" place="5" resultid="28466" />
                    <RANKING order="6" place="6" resultid="29258" />
                    <RANKING order="7" place="7" resultid="28842" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="12239" agemax="49" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="28849" />
                    <RANKING order="2" place="2" resultid="28225" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1195" agemax="98" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="29357" />
                    <RANKING order="2" place="2" resultid="28115" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="24851" daytime="14:55" gender="F" number="31" order="18" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="SURFACE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="24859" agemax="11" agemin="1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="29272" />
                    <RANKING order="2" place="2" resultid="28493" />
                    <RANKING order="3" place="3" resultid="29284" />
                    <RANKING order="4" place="4" resultid="28245" />
                    <RANKING order="5" place="5" resultid="29322" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="24852" agemax="13" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="29290" />
                    <RANKING order="2" place="2" resultid="28768" />
                    <RANKING order="3" place="3" resultid="29145" />
                    <RANKING order="4" place="4" resultid="28266" />
                    <RANKING order="5" place="5" resultid="29315" />
                    <RANKING order="6" place="-1" resultid="29278" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="24853" agemax="15" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="28712" />
                    <RANKING order="2" place="2" resultid="28717" />
                    <RANKING order="3" place="3" resultid="28503" />
                    <RANKING order="4" place="4" resultid="28514" />
                    <RANKING order="5" place="4" resultid="29238" />
                    <RANKING order="6" place="6" resultid="28259" />
                    <RANKING order="7" place="7" resultid="28508" />
                    <RANKING order="8" place="8" resultid="28498" />
                    <RANKING order="9" place="9" resultid="28471" />
                    <RANKING order="10" place="10" resultid="29308" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="24854" agemax="17" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="29223" />
                    <RANKING order="2" place="2" resultid="29188" />
                    <RANKING order="3" place="-1" resultid="29099" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="24855" agemax="34" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="28941" />
                    <RANKING order="2" place="2" resultid="28290" />
                    <RANKING order="3" place="3" resultid="28140" />
                    <RANKING order="4" place="-1" resultid="29296" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="24856" agemax="49" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="29327" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="24857" agemax="98" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="28441" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="24862" daytime="15:20" gender="M" number="32" order="19" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="SURFACE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="24863" agemax="11" agemin="1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="29103" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="24864" agemax="13" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="28529" />
                    <RANKING order="2" place="2" resultid="28766" />
                    <RANKING order="3" place="3" resultid="29341" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="24865" agemax="15" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="28701" />
                    <RANKING order="2" place="2" resultid="29228" />
                    <RANKING order="3" place="3" resultid="29116" />
                    <RANKING order="4" place="-1" resultid="29243" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="24866" agemax="17" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="28855" />
                    <RANKING order="2" place="2" resultid="28695" />
                    <RANKING order="3" place="3" resultid="29253" />
                    <RANKING order="4" place="4" resultid="28534" />
                    <RANKING order="5" place="5" resultid="29109" />
                    <RANKING order="6" place="6" resultid="29196" />
                    <RANKING order="7" place="7" resultid="28217" />
                    <RANKING order="8" place="-1" resultid="29204" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="24867" agemax="34" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="28689" />
                    <RANKING order="2" place="2" resultid="28176" />
                    <RANKING order="3" place="3" resultid="29209" />
                    <RANKING order="4" place="4" resultid="28170" />
                    <RANKING order="5" place="5" resultid="28124" />
                    <RANKING order="6" place="6" resultid="28196" />
                    <RANKING order="7" place="7" resultid="28183" />
                    <RANKING order="8" place="8" resultid="29374" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="24868" agemax="49" agemin="35" />
                <AGEGROUP agegroupid="24869" agemax="98" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="29358" />
                    <RANKING order="2" place="2" resultid="29334" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="1217" daytime="15:45" gender="F" number="33" order="22" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="4" stroke="SURFACE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1218" agemax="11" agemin="1" calculate="TOTAL" />
                <AGEGROUP agegroupid="1219" agemax="13" agemin="12" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="29380" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1220" agemax="15" agemin="14" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="29395" />
                    <RANKING order="2" place="2" resultid="29494" />
                    <RANKING order="3" place="3" resultid="28541" />
                    <RANKING order="4" place="4" resultid="28297" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1221" agemax="17" agemin="16" calculate="TOTAL" />
                <AGEGROUP agegroupid="1222" agemax="34" agemin="18" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="29378" />
                    <RANKING order="2" place="2" resultid="29387" />
                    <RANKING order="3" place="3" resultid="29493" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="12241" agemax="49" agemin="35" calculate="TOTAL" />
                <AGEGROUP agegroupid="1223" agemax="98" agemin="50" calculate="TOTAL" />
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="24873" daytime="15:55" gender="M" number="34" order="23" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="4" stroke="SURFACE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="24874" agemax="11" agemin="1" calculate="TOTAL" />
                <AGEGROUP agegroupid="24875" agemax="13" agemin="12" calculate="TOTAL" />
                <AGEGROUP agegroupid="24876" agemax="15" agemin="14" calculate="TOTAL" />
                <AGEGROUP agegroupid="24877" agemax="17" agemin="16" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="29123" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="24878" agemax="34" agemin="18" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="29396" />
                    <RANKING order="2" place="2" resultid="29484" />
                    <RANKING order="3" place="-1" resultid="29376" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="24879" agemax="49" agemin="35" calculate="TOTAL" />
                <AGEGROUP agegroupid="24880" agemax="98" agemin="50" calculate="TOTAL" />
              </AGEGROUPS>
            </EVENT>
          </EVENTS>
          <JUDGES>
            <JUDGE officialid="2149" remarks="ok" />
            <JUDGE officialid="21300" remarks="ok" />
            <JUDGE officialid="24070" remarks="ok" />
            <JUDGE officialid="28781" remarks="ok" />
            <JUDGE officialid="1520" remarks="ok" />
            <JUDGE officialid="25526" remarks="ok" />
            <JUDGE officialid="6661" remarks="ok" />
            <JUDGE officialid="1510" remarks="ok" />
            <JUDGE officialid="28777" remarks="ok" />
            <JUDGE officialid="2140" remarks="ok" />
            <JUDGE officialid="21335" remarks="ok" />
            <JUDGE officialid="26602" remarks="ok" />
            <JUDGE officialid="1538" remarks="ok" />
            <JUDGE number="101" officialid="4863" remarks="ok" />
            <JUDGE number="102" officialid="29471" remarks="ok" />
            <JUDGE number="103" officialid="25528" remarks="ok" />
            <JUDGE number="104" officialid="23071" remarks="ok" />
            <JUDGE number="204" officialid="28487" remarks="ok" />
            <JUDGE number="105" officialid="2148" remarks="ok" />
            <JUDGE number="106" officialid="5128" remarks="ok" />
            <JUDGE number="107" officialid="25527" remarks="ok" />
            <JUDGE number="108" officialid="27674" remarks="ok" />
            <JUDGE number="1" officialid="6383" remarks="OCEANUS" />
            <JUDGE number="2" officialid="3072" remarks="Orka &apos;97" />
            <JUDGE number="3" officialid="4401" remarks="OSV Delphis en Emese" />
            <JUDGE number="4" officialid="3074" remarks="OWT PONTOS" />
            <JUDGE number="5" officialid="3073" remarks="VZ Utrecht" />
            <JUDGE number="6" officialid="27676" remarks="Waves" />
            <JUDGE number="7" officialid="1536" remarks="MonoVinzz" />
            <JUDGE number="8" officialid="24198" remarks="DJK-VfR Muhlheim" />
            <JUDGE number="9" officialid="24196" remarks="TC Heilbronn" />
            <JUDGE number="10" officialid="24200" remarks="CS Gravenchon" />
            <JUDGE number="11" officialid="28804" remarks="SC DHfK Leipzig" />
            <JUDGE number="12" officialid="28804" remarks="TC Delitzsch" />
            <JUDGE number="13" officialid="28803" remarks="1. Chemnitz TVeV" />
            <JUDGE number="14" officialid="29436" remarks="Swiss Team" />
            <JUDGE number="15" officialid="27686" remarks="TC Nemo Plauen" />
            <JUDGE number="16" officialid="27807" remarks="PF NAP Aix" />
            <JUDGE number="17" officialid="28824" remarks="CSA Kremlin Bicetre" />
            <JUDGE number="18" officialid="24572" remarks="Tours NAP" />
            <JUDGE number="19" officialid="24482" remarks="Club Ciotaden NP" />
            <JUDGE number="20" officialid="27826" remarks="CPB NAP" />
            <JUDGE number="21" officialid="27683" remarks="Binger TSCeV" />
            <JUDGE number="22" officialid="24196" remarks="TC Harz" />
            <JUDGE number="23" officialid="24569" remarks="TC fez Berlin" />
            <JUDGE number="24" officialid="29179" remarks="LGM" />
            <JUDGE number="25" officialid="24573" remarks="Nautilus" />
            <JUDGE number="26" officialid="24795" remarks="Aq-Nivelles" />
          </JUDGES>
        </SESSION>
      </SESSIONS>
      <CLUBS>
        <CLUB type="CLUB" code="TCFB" nation="GER" clubid="22411" name="TC fez Berlin">
          <ATHLETES>
            <ATHLETE firstname="Rufus" lastname="Patge" birthdate="2006-05-15" gender="M" nation="GER" athleteid="29248">
              <RESULTS>
                <RESULT eventid="26746" points="952" reactiontime="+111" swimtime="00:08:14.58" resultid="29249" entrytime="00:08:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.02" />
                    <SPLIT distance="100" swimtime="00:00:56.63" />
                    <SPLIT distance="150" swimtime="00:01:27.16" />
                    <SPLIT distance="200" swimtime="00:01:58.06" />
                    <SPLIT distance="250" swimtime="00:02:28.47" />
                    <SPLIT distance="300" swimtime="00:03:00.00" />
                    <SPLIT distance="350" swimtime="00:03:31.39" />
                    <SPLIT distance="400" swimtime="00:04:02.37" />
                    <SPLIT distance="450" swimtime="00:04:35.21" />
                    <SPLIT distance="500" swimtime="00:05:06.57" />
                    <SPLIT distance="550" swimtime="00:05:38.14" />
                    <SPLIT distance="600" swimtime="00:06:09.81" />
                    <SPLIT distance="650" swimtime="00:06:41.91" />
                    <SPLIT distance="700" swimtime="00:07:13.32" />
                    <SPLIT distance="750" swimtime="00:07:44.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="7264" points="770" reactiontime="+90" swimtime="00:03:49.05" resultid="29250" entrytime="00:04:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:24.70" />
                    <SPLIT distance="100" swimtime="00:00:52.17" />
                    <SPLIT distance="150" swimtime="00:01:21.13" />
                    <SPLIT distance="200" swimtime="00:01:51.21" />
                    <SPLIT distance="250" swimtime="00:02:20.95" />
                    <SPLIT distance="300" swimtime="00:02:51.47" />
                    <SPLIT distance="350" swimtime="00:03:20.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="16574" points="724" reactiontime="+96" swimtime="00:08:15.99" resultid="29251" entrytime="00:08:01.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.82" />
                    <SPLIT distance="100" swimtime="00:00:57.90" />
                    <SPLIT distance="150" swimtime="00:01:28.07" />
                    <SPLIT distance="200" swimtime="00:01:59.00" />
                    <SPLIT distance="250" swimtime="00:02:30.27" />
                    <SPLIT distance="300" swimtime="00:03:01.82" />
                    <SPLIT distance="350" swimtime="00:03:33.96" />
                    <SPLIT distance="400" swimtime="00:04:06.30" />
                    <SPLIT distance="450" swimtime="00:04:38.04" />
                    <SPLIT distance="500" swimtime="00:05:08.64" />
                    <SPLIT distance="550" swimtime="00:05:40.14" />
                    <SPLIT distance="600" swimtime="00:06:12.53" />
                    <SPLIT distance="650" swimtime="00:06:43.17" />
                    <SPLIT distance="700" swimtime="00:07:14.55" />
                    <SPLIT distance="750" swimtime="00:07:45.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1203" points="684" reactiontime="+81" swimtime="00:04:29.78" resultid="29252" entrytime="00:04:48.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.32" />
                    <SPLIT distance="100" swimtime="00:01:03.23" />
                    <SPLIT distance="150" swimtime="00:01:36.85" />
                    <SPLIT distance="200" swimtime="00:02:12.19" />
                    <SPLIT distance="250" swimtime="00:02:47.65" />
                    <SPLIT distance="300" swimtime="00:03:22.59" />
                    <SPLIT distance="350" swimtime="00:03:57.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="24862" points="893" reactiontime="+89" swimtime="00:01:46.46" resultid="29253" entrytime="00:01:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:24.34" />
                    <SPLIT distance="100" swimtime="00:00:50.79" />
                    <SPLIT distance="150" swimtime="00:01:19.74" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Johanna" lastname="Schikora" birthdate="2002-01-06" gender="F" nation="GER" athleteid="29259">
              <RESULTS>
                <RESULT eventid="1093" points="1325" reactiontime="+101" swimtime="00:13:42.98" resultid="29260" entrytime="00:13:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.98" />
                    <SPLIT distance="100" swimtime="00:00:54.23" />
                    <SPLIT distance="150" swimtime="00:01:20.62" />
                    <SPLIT distance="200" swimtime="00:01:47.18" />
                    <SPLIT distance="250" swimtime="00:02:14.45" />
                    <SPLIT distance="300" swimtime="00:02:42.03" />
                    <SPLIT distance="350" swimtime="00:03:09.53" />
                    <SPLIT distance="400" swimtime="00:03:37.30" />
                    <SPLIT distance="450" swimtime="00:04:05.15" />
                    <SPLIT distance="500" swimtime="00:04:33.04" />
                    <SPLIT distance="550" swimtime="00:04:59.87" />
                    <SPLIT distance="600" swimtime="00:05:26.75" />
                    <SPLIT distance="650" swimtime="00:05:54.78" />
                    <SPLIT distance="700" swimtime="00:06:22.70" />
                    <SPLIT distance="750" swimtime="00:06:50.34" />
                    <SPLIT distance="800" swimtime="00:07:18.23" />
                    <SPLIT distance="850" swimtime="00:07:46.21" />
                    <SPLIT distance="900" swimtime="00:08:13.94" />
                    <SPLIT distance="950" swimtime="00:08:41.63" />
                    <SPLIT distance="1000" swimtime="00:09:09.48" />
                    <SPLIT distance="1050" swimtime="00:09:37.08" />
                    <SPLIT distance="1100" swimtime="00:10:04.89" />
                    <SPLIT distance="1150" swimtime="00:10:32.50" />
                    <SPLIT distance="1200" swimtime="00:11:00.03" />
                    <SPLIT distance="1250" swimtime="00:11:27.84" />
                    <SPLIT distance="1300" swimtime="00:11:55.83" />
                    <SPLIT distance="1350" swimtime="00:12:23.77" />
                    <SPLIT distance="1400" swimtime="00:12:51.18" />
                    <SPLIT distance="1450" swimtime="00:13:17.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1158" points="1277" reactiontime="+99" swimtime="00:07:11.59" resultid="29261" entrytime="00:06:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.05" />
                    <SPLIT distance="100" swimtime="00:00:54.08" />
                    <SPLIT distance="150" swimtime="00:01:20.75" />
                    <SPLIT distance="200" swimtime="00:01:47.12" />
                    <SPLIT distance="250" swimtime="00:02:14.38" />
                    <SPLIT distance="300" swimtime="00:02:41.68" />
                    <SPLIT distance="350" swimtime="00:03:09.15" />
                    <SPLIT distance="400" swimtime="00:03:36.68" />
                    <SPLIT distance="450" swimtime="00:04:04.18" />
                    <SPLIT distance="500" swimtime="00:04:31.48" />
                    <SPLIT distance="550" swimtime="00:04:58.48" />
                    <SPLIT distance="600" swimtime="00:05:25.58" />
                    <SPLIT distance="650" swimtime="00:05:53.09" />
                    <SPLIT distance="700" swimtime="00:06:20.30" />
                    <SPLIT distance="750" swimtime="00:06:46.73" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rèmy" lastname="Lebeau" birthdate="2002-05-28" gender="M" nation="FRA" athleteid="29254">
              <RESULTS>
                <RESULT eventid="26746" points="943" reactiontime="+124" swimtime="00:06:54.54" resultid="29255" entrytime="00:06:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:21.88" />
                    <SPLIT distance="100" swimtime="00:00:46.55" />
                    <SPLIT distance="150" swimtime="00:01:11.92" />
                    <SPLIT distance="200" swimtime="00:01:36.98" />
                    <SPLIT distance="250" swimtime="00:02:02.05" />
                    <SPLIT distance="300" swimtime="00:02:27.34" />
                    <SPLIT distance="350" swimtime="00:02:52.40" />
                    <SPLIT distance="400" swimtime="00:03:17.76" />
                    <SPLIT distance="450" swimtime="00:03:43.80" />
                    <SPLIT distance="500" swimtime="00:04:09.42" />
                    <SPLIT distance="550" swimtime="00:04:35.92" />
                    <SPLIT distance="600" swimtime="00:05:02.80" />
                    <SPLIT distance="650" swimtime="00:05:30.41" />
                    <SPLIT distance="700" swimtime="00:05:59.32" />
                    <SPLIT distance="750" swimtime="00:06:27.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1114" points="1168" reactiontime="+123" swimtime="00:03:03.09" resultid="29256" entrytime="00:03:00.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:21.20" />
                    <SPLIT distance="100" swimtime="00:00:43.90" />
                    <SPLIT distance="150" swimtime="00:01:07.09" />
                    <SPLIT distance="200" swimtime="00:01:30.81" />
                    <SPLIT distance="250" swimtime="00:01:54.74" />
                    <SPLIT distance="300" swimtime="00:02:18.06" />
                    <SPLIT distance="350" swimtime="00:02:40.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="16574" points="861" reactiontime="+96" swimtime="00:07:13.85" resultid="29257" entrytime="00:06:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:22.99" />
                    <SPLIT distance="100" swimtime="00:00:48.13" />
                    <SPLIT distance="150" swimtime="00:01:14.37" />
                    <SPLIT distance="200" swimtime="00:01:41.27" />
                    <SPLIT distance="250" swimtime="00:02:08.63" />
                    <SPLIT distance="300" swimtime="00:02:35.86" />
                    <SPLIT distance="350" swimtime="00:03:03.36" />
                    <SPLIT distance="400" swimtime="00:03:30.97" />
                    <SPLIT distance="450" swimtime="00:03:58.60" />
                    <SPLIT distance="500" swimtime="00:04:26.65" />
                    <SPLIT distance="550" swimtime="00:04:54.58" />
                    <SPLIT distance="600" swimtime="00:05:22.56" />
                    <SPLIT distance="650" swimtime="00:05:51.03" />
                    <SPLIT distance="700" swimtime="00:06:19.40" />
                    <SPLIT distance="750" swimtime="00:06:47.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1190" points="540" reactiontime="+117" swimtime="00:00:44.87" resultid="29258" entrytime="00:00:38.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:22.76" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <OFFICIALS>
            <OFFICIAL officialid="24569" firstname="Volko" gender="M" grade="Team Captain" lastname="Kucher" nation="GER" />
          </OFFICIALS>
        </CLUB>
        <CLUB type="CLUB" code="RIESA/DRES" clubid="22889" name="RIESA/DRESDEN" />
        <CLUB type="CLUB" code="ORKA&apos;97" nation="NED" clubid="16851" name="Orka &apos;97">
          <ATHLETES>
            <ATHLETE firstname="Rianne" lastname="Smit" birthdate="1997-10-29" gender="F" nation="NED" license="9024377" athleteid="28132">
              <RESULTS>
                <RESULT eventid="1053" points="416" reactiontime="+85" swimtime="00:00:26.73" resultid="28133" entrytime="00:00:27.55" entrycourse="LCM" />
                <RESULT eventid="7254" points="502" reactiontime="+82" swimtime="00:02:19.02" resultid="28134" entrytime="00:02:28.83" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.30" />
                    <SPLIT distance="100" swimtime="00:01:05.91" />
                    <SPLIT distance="150" swimtime="00:01:42.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1120" points="594" reactiontime="+82" swimtime="00:00:27.74" resultid="28135" entrytime="00:00:29.62" entrycourse="LCM" />
                <RESULT eventid="7278" points="357" reactiontime="+102" swimtime="00:05:15.79" resultid="28136" entrytime="00:05:10.02" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.48" />
                    <SPLIT distance="100" swimtime="00:01:12.11" />
                    <SPLIT distance="150" swimtime="00:01:52.36" />
                    <SPLIT distance="200" swimtime="00:02:33.13" />
                    <SPLIT distance="250" swimtime="00:03:14.94" />
                    <SPLIT distance="300" swimtime="00:03:56.63" />
                    <SPLIT distance="350" swimtime="00:04:38.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1168" points="572" reactiontime="+82" swimtime="00:01:01.19" resultid="28137" entrytime="00:01:03.32" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="7287" points="406" reactiontime="+95" swimtime="00:01:01.97" resultid="28138" entrytime="00:01:02.49" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1196" points="598" reactiontime="+86" swimtime="00:05:13.30" resultid="28139" entrytime="00:05:24.41" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.69" />
                    <SPLIT distance="100" swimtime="00:01:15.42" />
                    <SPLIT distance="150" swimtime="00:01:55.48" />
                    <SPLIT distance="200" swimtime="00:02:36.52" />
                    <SPLIT distance="250" swimtime="00:03:17.01" />
                    <SPLIT distance="300" swimtime="00:03:58.35" />
                    <SPLIT distance="350" swimtime="00:04:37.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="24851" points="330" reactiontime="+100" swimtime="00:02:26.57" resultid="28140">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.29" />
                    <SPLIT distance="100" swimtime="00:01:08.85" />
                    <SPLIT distance="150" swimtime="00:01:49.27" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Tara" lastname="Graafland" birthdate="2001-01-16" gender="F" nation="NED" license="9035812" athleteid="28125">
              <RESULTS>
                <RESULT eventid="1147" points="465" reactiontime="+118" swimtime="00:00:24.33" resultid="28126" entrytime="00:00:24.23" entrycourse="LCM" />
                <RESULT eventid="1168" points="611" reactiontime="+103" swimtime="00:00:59.86" resultid="28127" entrytime="00:01:01.45" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="7287" points="490" reactiontime="+100" swimtime="00:00:58.23" resultid="28128" entrytime="00:00:58.93" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.19" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Eva" lastname="Moolenkamp" birthdate="2008-06-01" gender="F" nation="NED" license="9265760" athleteid="28129">
              <RESULTS>
                <RESULT eventid="1053" points="380" reactiontime="+94" swimtime="00:00:29.57" resultid="28130" entrytime="00:00:29.71" entrycourse="LCM" />
                <RESULT eventid="1120" points="502" reactiontime="+98" swimtime="00:00:31.24" resultid="28131" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Peter" lastname="Blanker" birthdate="1972-04-23" gender="M" nation="NED" license="35291" athleteid="28110">
              <RESULTS>
                <RESULT eventid="1079" points="548" reactiontime="+126" swimtime="00:00:25.97" resultid="28111" entrytime="00:00:28.14" entrycourse="LCM" />
                <RESULT eventid="7271" points="762" reactiontime="+102" swimtime="00:02:08.69" resultid="28112">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.42" />
                    <SPLIT distance="100" swimtime="00:01:00.29" />
                    <SPLIT distance="150" swimtime="00:01:34.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1114" points="519" reactiontime="+143" swimtime="00:05:09.10" resultid="28113" entrytime="00:05:12.25" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.31" />
                    <SPLIT distance="100" swimtime="00:01:09.87" />
                    <SPLIT distance="150" swimtime="00:01:49.07" />
                    <SPLIT distance="200" swimtime="00:02:29.80" />
                    <SPLIT distance="250" swimtime="00:03:10.20" />
                    <SPLIT distance="300" swimtime="00:03:51.50" />
                    <SPLIT distance="350" swimtime="00:04:32.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="16574" points="565" reactiontime="+110" swimtime="00:10:02.92" resultid="28114">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.43" />
                    <SPLIT distance="100" swimtime="00:01:07.05" />
                    <SPLIT distance="150" swimtime="00:01:45.00" />
                    <SPLIT distance="200" swimtime="00:02:24.08" />
                    <SPLIT distance="250" swimtime="00:03:03.00" />
                    <SPLIT distance="300" swimtime="00:03:41.96" />
                    <SPLIT distance="350" swimtime="00:04:21.23" />
                    <SPLIT distance="400" swimtime="00:05:00.64" />
                    <SPLIT distance="450" swimtime="00:05:39.63" />
                    <SPLIT distance="500" swimtime="00:06:18.84" />
                    <SPLIT distance="550" swimtime="00:06:57.45" />
                    <SPLIT distance="600" swimtime="00:07:36.41" />
                    <SPLIT distance="650" swimtime="00:08:14.90" />
                    <SPLIT distance="700" swimtime="00:08:53.69" />
                    <SPLIT distance="750" swimtime="00:09:29.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1190" points="555" reactiontime="+120" swimtime="00:00:57.70" resultid="28115" entrytime="00:01:00.52" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.47" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Roelant" lastname="Cornelissen" birthdate="1991-10-08" gender="M" nation="NED" license="9259164" athleteid="28116">
              <RESULTS>
                <RESULT eventid="1079" points="432" reactiontime="+97" swimtime="00:00:22.41" resultid="28117" entrytime="00:00:22.08" entrycourse="LCM" />
                <RESULT eventid="7271" points="796" reactiontime="+87" swimtime="00:01:57.54" resultid="28118" entrytime="00:01:55.93" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.84" />
                    <SPLIT distance="100" swimtime="00:00:56.27" />
                    <SPLIT distance="150" swimtime="00:01:27.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1127" points="656" reactiontime="+86" swimtime="00:00:23.24" resultid="28119" entrytime="00:00:23.77" entrycourse="LCM" />
                <RESULT eventid="7264" points="442" reactiontime="+107" swimtime="00:04:17.96" resultid="28120" entrytime="00:04:20.31" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.08" />
                    <SPLIT distance="100" swimtime="00:00:59.82" />
                    <SPLIT distance="150" swimtime="00:01:32.11" />
                    <SPLIT distance="200" swimtime="00:02:05.23" />
                    <SPLIT distance="250" swimtime="00:02:38.70" />
                    <SPLIT distance="300" swimtime="00:03:13.05" />
                    <SPLIT distance="350" swimtime="00:03:46.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1153" points="576" reactiontime="+107" swimtime="00:00:19.00" resultid="28121" entrytime="00:00:20.12" entrycourse="LCM" />
                <RESULT eventid="1175" points="720" reactiontime="+90" swimtime="00:00:51.49" resultid="28122">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:24.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1203" points="600" reactiontime="+97" swimtime="00:04:31.33" resultid="28123" entrytime="00:04:58.78" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.89" />
                    <SPLIT distance="100" swimtime="00:01:04.02" />
                    <SPLIT distance="150" swimtime="00:01:39.18" />
                    <SPLIT distance="200" swimtime="00:02:14.05" />
                    <SPLIT distance="250" swimtime="00:02:49.35" />
                    <SPLIT distance="300" swimtime="00:03:24.09" />
                    <SPLIT distance="350" swimtime="00:03:59.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="24862" points="525" reactiontime="+102" swimtime="00:01:53.93" resultid="28124">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.00" />
                    <SPLIT distance="100" swimtime="00:00:52.89" />
                    <SPLIT distance="150" swimtime="00:01:23.87" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <OFFICIALS>
            <OFFICIAL officialid="7491" firstname="Annette" gender="F" grade="Kamprechter" lastname="Groot" nameprefix="de" nation="NED" />
            <OFFICIAL officialid="7618" firstname="dochter" gender="F" grade="briefloper" lastname="Hove" nameprefix="ten" nation="NED" />
            <OFFICIAL officialid="6380" firstname="Michael" grade="gastheer DOV Botlek" lastname="Ruisch" nation="NED" />
            <OFFICIAL officialid="4866" firstname="Adri" gender="M" grade="Hulp secretariaat" lastname="Broersen" nation="NED" />
            <OFFICIAL officialid="7842" firstname="Marly" gender="F" grade="kamprechter" lastname="Smit" nation="NED" />
            <OFFICIAL officialid="24074" firstname="Jeoffry" gender="M" grade="Tijdwaarnemer" lastname="Esch" nameprefix="van" nation="NED" />
            <OFFICIAL officialid="1527" firstname="Jeoffry" gender="M" grade="Lijnrechter" lastname="Esch" nameprefix="van" nation="NED" />
            <OFFICIAL officialid="4850" firstname="Angelo" gender="M" grade="gastheer DOV Botlek" lastname="Eikmans" nation="NED" />
            <OFFICIAL officialid="4870" firstname="Jolanda" gender="F" grade="Speaker" lastname="Doeselaar" nameprefix="van" nation="NED" />
            <OFFICIAL officialid="3072" firstname="Peter" grade="Ploegleider" lastname="Blanker" nation="NED" />
            <OFFICIAL officialid="23170" firstname="Gerard" gender="M" grade="Speaker" lastname="Veurink" nation="NED" />
            <OFFICIAL officialid="4851" firstname="Gerard" gender="M" grade="Starter" lastname="Veurink" nation="NED" />
            <OFFICIAL officialid="2141" firstname="Johan" gender="M" grade="EHB(D)O" lastname="Herwijnen" nation="NED" />
            <OFFICIAL officialid="6372" firstname="Annet" gender="F" grade="Kamprechter" lastname="Groot" nameprefix="de" nation="NED" />
            <OFFICIAL officialid="24070" firstname="Peter" gender="M" grade="Wedstrijd indeling" lastname="Blanker" nation="NED" />
          </OFFICIALS>
        </CLUB>
        <CLUB type="CLUB" code="PCD" nation="FRA" clubid="21969" name="Plongée Club de Douai" />
        <CLUB type="CLUB" code="TMP" nation="FRA" clubid="27620" name="Toulouse Métropole Palmes">
          <OFFICIALS>
            <OFFICIAL officialid="27690" firstname="Delphine" gender="F" grade="Team Captain" lastname="Dujardin" nation="FRA" />
          </OFFICIALS>
        </CLUB>
        <CLUB type="CLUB" code="DSF" nation="DEN" clubid="22500" name="Dansk Sportsdykker Forbund">
          <OFFICIALS>
            <OFFICIAL officialid="24203" firstname="Kenneth" gender="M" grade="Team Captain" lastname="Aaberg" nation="DEN" />
          </OFFICIALS>
        </CLUB>
        <CLUB type="CLUB" code="DAW" nation="NED" clubid="18181" name="DAW Alkmaar">
          <OFFICIALS>
            <OFFICIAL officialid="1520" firstname="Leo" grade="Vz. Kamprechter" lastname="Bol" nation="NED" />
            <OFFICIAL officialid="1511" firstname="Niek" gender="M" grade="Tijdwaarnemer" lastname="Kloots" nation="NED" />
            <OFFICIAL officialid="1521" firstname="Karel" grade="Tijdwaarnemer" lastname="Bol" nation="NED" />
          </OFFICIALS>
        </CLUB>
        <CLUB type="CLUB" code="BELGIUM" clubid="24809" name="Belgium" />
        <CLUB type="CLUB" code="SCRF" nation="GER" clubid="22873" name="SC Riesa Finswimming" />
        <CLUB type="CLUB" code="ZVH" nation="NED" clubid="20111" name="ZV Hoogland">
          <OFFICIALS>
            <OFFICIAL officialid="21320" firstname="Ada" gender="F" grade="Tijdwaarnemer" lastname="Smit" nameprefix="de" nation="NED" />
            <OFFICIAL officialid="25526" firstname="Ada" gender="F" grade="( VZ) Kamprechter" lastname="Smit" nameprefix="de" nation="NED" />
            <OFFICIAL officialid="23287" firstname="Diego" gender="M" grade="Ploegleider" lastname="Quintero" nation="NED" />
          </OFFICIALS>
        </CLUB>
        <CLUB type="CLUB" code="TSCB" nation="GER" clubid="22870" name="Berliner TSC" />
        <CLUB type="CLUB" code="OSV DELPHI" nation="NED" clubid="23286" name="OSV Delphis">
          <ATHLETES>
            <ATHLETE firstname="Nerena" lastname="Vuuren" birthdate="2002-06-28" gender="F" nameprefix="van" nation="NED" license="9010785" athleteid="28141">
              <RESULTS>
                <RESULT eventid="1093" points="378" reactiontime="+120" swimtime="00:20:49.35" resultid="28142" entrytime="00:20:43.92" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.78" />
                    <SPLIT distance="100" swimtime="00:01:10.46" />
                    <SPLIT distance="150" swimtime="00:01:51.02" />
                    <SPLIT distance="200" swimtime="00:02:32.77" />
                    <SPLIT distance="250" swimtime="00:03:14.07" />
                    <SPLIT distance="300" swimtime="00:03:56.01" />
                    <SPLIT distance="350" swimtime="00:04:38.16" />
                    <SPLIT distance="400" swimtime="00:05:20.66" />
                    <SPLIT distance="450" swimtime="00:06:02.64" />
                    <SPLIT distance="500" swimtime="00:06:44.66" />
                    <SPLIT distance="550" swimtime="00:07:26.77" />
                    <SPLIT distance="600" swimtime="00:08:08.36" />
                    <SPLIT distance="650" swimtime="00:08:51.23" />
                    <SPLIT distance="700" swimtime="00:09:33.08" />
                    <SPLIT distance="750" swimtime="00:10:15.09" />
                    <SPLIT distance="800" swimtime="00:10:57.03" />
                    <SPLIT distance="850" swimtime="00:11:39.83" />
                    <SPLIT distance="900" swimtime="00:12:23.63" />
                    <SPLIT distance="950" swimtime="00:13:05.72" />
                    <SPLIT distance="1000" swimtime="00:13:48.46" />
                    <SPLIT distance="1050" swimtime="00:14:32.12" />
                    <SPLIT distance="1100" swimtime="00:15:15.34" />
                    <SPLIT distance="1150" swimtime="00:15:57.73" />
                    <SPLIT distance="1200" swimtime="00:16:42.02" />
                    <SPLIT distance="1250" swimtime="00:17:24.25" />
                    <SPLIT distance="1300" swimtime="00:18:07.52" />
                    <SPLIT distance="1350" swimtime="00:18:49.68" />
                    <SPLIT distance="1400" swimtime="00:19:31.29" />
                    <SPLIT distance="1450" swimtime="00:20:11.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="7254" points="402" reactiontime="+108" swimtime="00:02:29.73" resultid="28143" entrytime="00:02:20.51" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.52" />
                    <SPLIT distance="100" swimtime="00:01:08.81" />
                    <SPLIT distance="150" swimtime="00:01:50.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1120" points="573" reactiontime="+98" swimtime="00:00:28.08" resultid="28144" entrytime="00:00:28.37" entrycourse="LCM" />
                <RESULT eventid="1105" points="257" reactiontime="+143" swimtime="00:05:49.63" resultid="28145" entrytime="00:05:39.51" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.23" />
                    <SPLIT distance="100" swimtime="00:01:22.65" />
                    <SPLIT distance="150" swimtime="00:02:08.50" />
                    <SPLIT distance="200" swimtime="00:02:54.52" />
                    <SPLIT distance="250" swimtime="00:03:40.32" />
                    <SPLIT distance="300" swimtime="00:04:24.28" />
                    <SPLIT distance="350" swimtime="00:05:09.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1168" points="514" reactiontime="+104" swimtime="00:01:03.42" resultid="28146" entrytime="00:01:03.44" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1196" points="622" reactiontime="+111" swimtime="00:05:09.30" resultid="28147" entrytime="00:05:04.73" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.24" />
                    <SPLIT distance="100" swimtime="00:01:12.64" />
                    <SPLIT distance="150" swimtime="00:01:52.53" />
                    <SPLIT distance="200" swimtime="00:02:33.56" />
                    <SPLIT distance="250" swimtime="00:03:14.10" />
                    <SPLIT distance="300" swimtime="00:03:53.89" />
                    <SPLIT distance="350" swimtime="00:04:33.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1182" points="225" reactiontime="+136" swimtime="00:01:12.59" resultid="28148">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.05" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <OFFICIALS>
            <OFFICIAL officialid="29057" firstname="Marian" gender="F" grade="secretariaat (io)" lastname="Beukel" nameprefix="van den" nation="NED" />
            <OFFICIAL officialid="4401" firstname="Rene" gender="M" grade="Ploegleider" lastname="Vuuren" nameprefix="van" nation="NED" />
            <OFFICIAL officialid="7858" firstname="Marco" gender="M" grade="Lijnrechter" lastname="Beukel" nameprefix="van den" nation="NED" />
          </OFFICIALS>
        </CLUB>
        <CLUB type="CLUB" code="LGM" nation="BEL" clubid="22123" name="Liege Grivegnee Monopalme">
          <ATHLETES>
            <ATHLETE firstname="Aramé" lastname="Guevorkyan" birthdate="2007-01-01" gender="M" nation="BEL" license="55415" athleteid="29181">
              <RESULTS>
                <RESULT eventid="1079" reactiontime="+95" status="DSQ" swimtime="00:00:22.92" resultid="29193" entrytime="00:00:23.91" />
                <RESULT eventid="1127" points="615" reactiontime="+105" swimtime="00:00:26.58" resultid="29194" entrytime="00:00:25.00" />
                <RESULT eventid="7295" points="473" reactiontime="+98" swimtime="00:00:52.40" resultid="29195" entrytime="00:00:53.22">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:24.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="24862" points="557" reactiontime="+105" swimtime="00:02:04.60" resultid="29196" entrytime="00:02:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.26" />
                    <SPLIT distance="100" swimtime="00:00:59.66" />
                    <SPLIT distance="150" swimtime="00:01:32.92" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Sandra" lastname="Gallo" birthdate="2010-01-01" gender="F" nation="BEL" license="55416" athleteid="29180">
              <RESULTS>
                <RESULT eventid="1053" points="230" reactiontime="+126" swimtime="00:00:37.04" resultid="29189" entrytime="00:00:45.00" />
                <RESULT comment="A7 - Niet aangekomen met alle materialen, waarmee men vertrokken is" eventid="7254" reactiontime="+118" status="DSQ" swimtime="00:00:00.00" resultid="29190" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.52" />
                    <SPLIT distance="100" swimtime="00:01:28.45" />
                    <SPLIT distance="150" swimtime="00:02:27.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1168" points="426" reactiontime="+94" swimtime="00:01:18.55" resultid="29191" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="7287" points="218" reactiontime="+105" swimtime="00:01:23.34" resultid="29192" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.49" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Cassandra" lastname="Membert" birthdate="2006-01-01" gender="F" nation="BEL" license="55413" athleteid="29182">
              <RESULTS>
                <RESULT comment="A2 - Niet gestart" eventid="1053" status="DSQ" swimtime="00:00:00.00" resultid="29197" entrytime="00:00:32.52" />
                <RESULT eventid="7254" points="468" reactiontime="+92" swimtime="00:02:33.77" resultid="29198" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.66" />
                    <SPLIT distance="100" swimtime="00:01:11.78" />
                    <SPLIT distance="150" swimtime="00:01:54.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1168" points="491" reactiontime="+91" swimtime="00:01:07.42" resultid="29199" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="7287" points="346" reactiontime="+95" swimtime="00:01:05.85" resultid="29200" entrytime="00:01:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.40" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Cali" lastname="Poussart" birthdate="2007-01-01" gender="M" nation="BEL" license="55417" athleteid="29183">
              <RESULTS>
                <RESULT comment="A11 - Uitrusting voldoet niet aan de geldende eisen" eventid="1079" status="DSQ" swimtime="00:00:00.00" resultid="29201" entrytime="00:00:30.00" />
                <RESULT eventid="1175" points="630" reactiontime="+83" swimtime="00:00:58.54" resultid="29202" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.87" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="A3 - De aangegeven zwemwijze niet uitgevoerd (oa duiken)" eventid="7295" reactiontime="+105" status="DSQ" swimtime="00:00:00.00" resultid="29203" entrytime="00:01:02.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.77" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="A3 - De aangegeven zwemwijze niet uitgevoerd (oa duiken)" eventid="24862" reactiontime="+102" status="DSQ" swimtime="00:02:15.61" resultid="29204" entrytime="00:02:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.91" />
                    <SPLIT distance="100" swimtime="00:01:06.55" />
                    <SPLIT distance="150" swimtime="00:01:43.81" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Léonard" lastname="Alaimo" birthdate="1999-01-01" gender="M" nation="BEL" license="43895" athleteid="29184">
              <RESULTS>
                <RESULT eventid="1079" points="756" reactiontime="+94" swimtime="00:00:18.60" resultid="29205" entrytime="00:00:18.30" />
                <RESULT eventid="1127" points="733" reactiontime="+78" swimtime="00:00:22.40" resultid="29206" entrytime="00:00:21.50" />
                <RESULT eventid="1153" points="818" reactiontime="+92" swimtime="00:00:16.90" resultid="29207" entrytime="00:00:17.80" />
                <RESULT eventid="7295" points="858" reactiontime="+89" swimtime="00:00:41.48" resultid="29208" entrytime="00:00:40.06">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:19.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="24862" points="757" reactiontime="+90" swimtime="00:01:40.83" resultid="29209" entrytime="00:01:33.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:22.48" />
                    <SPLIT distance="100" swimtime="00:00:47.29" />
                    <SPLIT distance="150" swimtime="00:01:14.24" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Sarah" lastname="Gallo" birthdate="2007-01-01" gender="F" nation="BEL" license="48930" athleteid="29178">
              <RESULTS>
                <RESULT comment="A2 - Niet gestart" eventid="1053" status="DSQ" swimtime="00:00:00.00" resultid="29185" entrytime="00:00:31.97" />
                <RESULT eventid="7254" points="492" reactiontime="+101" swimtime="00:02:31.20" resultid="29186" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.58" />
                    <SPLIT distance="100" swimtime="00:01:09.14" />
                    <SPLIT distance="150" swimtime="00:01:51.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="7287" points="494" reactiontime="+111" swimtime="00:00:58.49" resultid="29187" entrytime="00:01:02.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="24851" points="428" reactiontime="+105" swimtime="00:02:17.02" resultid="29188" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.82" />
                    <SPLIT distance="100" swimtime="00:01:01.50" />
                    <SPLIT distance="150" swimtime="00:01:39.78" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="17" agemin="16" agetotalmax="-1" agetotalmin="-1" gender="X" name="LGM GB" number="1">
              <RESULTS>
                <RESULT eventid="1140" reactiontime="+93" swimtime="00:04:14.38" resultid="29210">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.52" />
                    <SPLIT distance="100" swimtime="00:00:57.28" />
                    <SPLIT distance="150" swimtime="00:01:31.19" />
                    <SPLIT distance="200" swimtime="00:02:07.35" />
                    <SPLIT distance="250" swimtime="00:02:35.93" />
                    <SPLIT distance="300" swimtime="00:03:07.49" />
                    <SPLIT distance="350" swimtime="00:03:39.11" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="29181" number="1" reactiontime="+93" />
                    <RELAYPOSITION athleteid="29182" number="2" reactiontime="+55" />
                    <RELAYPOSITION athleteid="29183" number="3" reactiontime="+16" />
                    <RELAYPOSITION athleteid="29178" number="4" reactiontime="+60" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
          <OFFICIALS>
            <OFFICIAL officialid="29179" firstname="Alaimo" gender="M" grade="Team Captain" lastname="Léonard" nation="BEL" />
            <OFFICIAL officialid="24480" firstname="Bruno" gender="M" grade="Team Captain" lastname="Dupont" nation="BEL" />
          </OFFICIALS>
        </CLUB>
        <CLUB type="CLUB" code="LIV FC" nation="INA" clubid="22876" name="LIV Finswimming club" shortname="LIV FC">
          <OFFICIALS>
            <OFFICIAL officialid="26646" firstname="Ciska" gender="F" grade="Team Captain" lastname="Herawati" nation="INA" />
          </OFFICIALS>
        </CLUB>
        <CLUB type="CLUB" code="NOB" nation="NED" clubid="17409" name="NOB">
          <ATHLETES>
            <ATHLETE firstname="Mahmoud" lastname="Hassan" birthdate="1991-08-17" gender="M" nation="NED" license="9265697" athleteid="28100">
              <RESULTS>
                <RESULT comment="A1 - Bewogen of te vroeg weg bij de start (geen tijd noteren)" eventid="7271" reactiontime="+78" status="DSQ" swimtime="00:01:49.13" resultid="28101" entrytime="00:01:54.47" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:24.81" />
                    <SPLIT distance="100" swimtime="00:00:51.84" />
                    <SPLIT distance="150" swimtime="00:01:20.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1127" points="739" reactiontime="+88" swimtime="00:00:22.34" resultid="28102" />
                <RESULT eventid="1175" points="863" reactiontime="+86" swimtime="00:00:48.48" resultid="28103" entrytime="00:00:50.63" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:23.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1203" points="797" reactiontime="+92" swimtime="00:04:06.81" resultid="28104" entrytime="00:04:36.45" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.49" />
                    <SPLIT distance="100" swimtime="00:00:56.14" />
                    <SPLIT distance="150" swimtime="00:01:27.21" />
                    <SPLIT distance="200" swimtime="00:01:59.08" />
                    <SPLIT distance="250" swimtime="00:02:31.22" />
                    <SPLIT distance="300" swimtime="00:03:03.89" />
                    <SPLIT distance="350" swimtime="00:03:36.57" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="34" agetotalmin="18" gender="M" name="NOB HA" number="1">
              <RESULTS>
                <RESULT eventid="26768" reactiontime="+85" swimtime="00:01:30.85" resultid="29473">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:22.30" />
                    <SPLIT distance="100" swimtime="00:00:44.49" />
                    <SPLIT distance="150" swimtime="00:01:04.77" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="28100" number="1" reactiontime="+85" />
                    <RELAYPOSITION athleteid="28116" number="2" reactiontime="+15" />
                    <RELAYPOSITION athleteid="29350" number="3" reactiontime="+47" />
                    <RELAYPOSITION athleteid="28110" number="4" reactiontime="+62" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="34" agetotalmin="18" gender="F" name="NOB DA" number="3">
              <RESULTS>
                <RESULT eventid="26758" reactiontime="+100" swimtime="00:01:48.56" resultid="29386">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.29" />
                    <SPLIT distance="100" swimtime="00:00:54.24" />
                    <SPLIT distance="150" swimtime="00:01:21.03" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="28252" number="1" reactiontime="+100" />
                    <RELAYPOSITION athleteid="28129" number="2" reactiontime="+2" />
                    <RELAYPOSITION athleteid="28282" number="3" reactiontime="+82" />
                    <RELAYPOSITION athleteid="28105" number="4" reactiontime="+65" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="34" agetotalmin="18" gender="F" name="NOB DA" number="3">
              <RESULTS>
                <RESULT eventid="1217" reactiontime="+119" swimtime="00:04:07.74" resultid="29387">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.30" />
                    <SPLIT distance="100" swimtime="00:00:58.00" />
                    <SPLIT distance="150" swimtime="00:01:28.11" />
                    <SPLIT distance="200" swimtime="00:02:02.20" />
                    <SPLIT distance="250" swimtime="00:02:32.68" />
                    <SPLIT distance="300" swimtime="00:03:07.91" />
                    <SPLIT distance="350" swimtime="00:03:37.11" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="28125" number="1" reactiontime="+119" />
                    <RELAYPOSITION athleteid="28132" number="2" reactiontime="+38" />
                    <RELAYPOSITION athleteid="28141" number="3" reactiontime="+71" />
                    <RELAYPOSITION athleteid="28105" number="4" reactiontime="+106" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="34" agemin="18" agetotalmax="-1" agetotalmin="-1" gender="X" name="NOB 3D1H BM">
              <RESULTS>
                <RESULT eventid="1140" reactiontime="+99" status="EXH" swimtime="00:04:13.76" resultid="29487" late="yes">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.45" />
                    <SPLIT distance="100" swimtime="00:01:10.31" />
                    <SPLIT distance="150" swimtime="00:01:41.73" />
                    <SPLIT distance="200" swimtime="00:02:16.49" />
                    <SPLIT distance="250" swimtime="00:02:44.05" />
                    <SPLIT distance="300" swimtime="00:03:14.65" />
                    <SPLIT distance="350" swimtime="00:03:43.42" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="28246" number="1" reactiontime="+99" />
                    <RELAYPOSITION athleteid="28282" number="2" reactiontime="+56" />
                    <RELAYPOSITION athleteid="28110" number="3" reactiontime="+66" />
                    <RELAYPOSITION athleteid="29285" number="4" reactiontime="+54" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="34" agemin="18" agetotalmax="-1" agetotalmin="-1" gender="X" name="NOB GA">
              <RESULTS>
                <RESULT eventid="1140" reactiontime="+84" swimtime="00:03:55.96" resultid="29488" late="yes">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.20" />
                    <SPLIT distance="100" swimtime="00:01:02.07" />
                    <SPLIT distance="150" swimtime="00:01:32.99" />
                    <SPLIT distance="200" swimtime="00:02:07.68" />
                    <SPLIT distance="250" swimtime="00:02:32.13" />
                    <SPLIT distance="300" swimtime="00:02:59.37" />
                    <SPLIT distance="350" swimtime="00:03:26.66" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="28132" number="1" reactiontime="+84" />
                    <RELAYPOSITION athleteid="28141" number="2" reactiontime="+71" />
                    <RELAYPOSITION athleteid="28116" number="3" reactiontime="+40" />
                    <RELAYPOSITION athleteid="28204" number="4" reactiontime="+46" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="34" agetotalmin="18" gender="X" name="NOB GA">
              <RESULTS>
                <RESULT eventid="1210" reactiontime="+106" swimtime="00:01:31.55" resultid="29492" late="yes">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:20.06" />
                    <SPLIT distance="100" swimtime="00:00:43.01" />
                    <SPLIT distance="150" swimtime="00:01:07.59" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="28116" number="1" reactiontime="+106" />
                    <RELAYPOSITION athleteid="29342" number="2" reactiontime="+39" />
                    <RELAYPOSITION athleteid="29368" number="3" reactiontime="+47" />
                    <RELAYPOSITION athleteid="29362" number="4" reactiontime="+31" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="34" agemin="18" agetotalmax="-1" agetotalmin="-1" gender="X" name="NOB GA PONTOS Mahmoud">
              <RESULTS>
                <RESULT eventid="1140" reactiontime="+89" swimtime="00:03:49.48" resultid="29490" late="yes">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:24.33" />
                    <SPLIT distance="100" swimtime="00:00:50.67" />
                    <SPLIT distance="150" swimtime="00:01:22.47" />
                    <SPLIT distance="200" swimtime="00:01:57.67" />
                    <SPLIT distance="250" swimtime="00:02:20.86" />
                    <SPLIT distance="300" swimtime="00:02:46.42" />
                    <SPLIT distance="350" swimtime="00:03:15.51" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="28231" number="1" reactiontime="+89" />
                    <RELAYPOSITION athleteid="28267" number="2" reactiontime="+19" />
                    <RELAYPOSITION athleteid="28100" number="3" reactiontime="+59" />
                    <RELAYPOSITION athleteid="28252" number="4" reactiontime="+48" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
          <OFFICIALS>
            <OFFICIAL officialid="4868" firstname="Alex" gender="M" grade="Briefloper" lastname="Diepen" nameprefix="van" nation="NED" />
            <OFFICIAL officialid="21329" firstname="Daniël" gender="M" grade="bestuurslid Sport" lastname="Bakel" nameprefix="van" nation="NED" />
            <OFFICIAL officialid="24072" firstname="Erik" gender="M" grade="Opening" lastname="Vessem" nameprefix="van" nation="NED" />
          </OFFICIALS>
        </CLUB>
        <CLUB type="CLUB" code="RELAY GER" nation="GER" clubid="24240" name="Relay Germany" shortname="RELAY GER">
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="34" agetotalmin="18" gender="M" name="Team Saxony HA" number="1">
              <RESULTS>
                <RESULT comment="B2 - Na start- en/of keerpunt meer dan 15 meter onder water gezwommen" eventid="26768" reactiontime="+82" status="DSQ" swimtime="00:01:13.88" resultid="29389" entrytime="00:01:13.01">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:18.11" />
                    <SPLIT distance="100" swimtime="00:00:37.91" />
                    <SPLIT distance="150" swimtime="00:00:56.95" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="28685" number="1" reactiontime="+82" status="DSQ" />
                    <RELAYPOSITION athleteid="28696" number="2" reactiontime="+52" status="DSQ" />
                    <RELAYPOSITION athleteid="28690" number="3" reactiontime="+56" status="DSQ" />
                    <RELAYPOSITION athleteid="27813" number="4" reactiontime="+16" status="DSQ" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="34" agetotalmin="18" gender="M" name="Team Saxony HA" number="1">
              <RESULTS>
                <RESULT eventid="24873" reactiontime="+81" swimtime="00:02:48.86" resultid="29396" entrytime="00:02:49.13">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:19.62" />
                    <SPLIT distance="100" swimtime="00:00:41.79" />
                    <SPLIT distance="150" swimtime="00:01:03.33" />
                    <SPLIT distance="200" swimtime="00:01:27.35" />
                    <SPLIT distance="250" swimtime="00:01:47.58" />
                    <SPLIT distance="300" swimtime="00:02:09.78" />
                    <SPLIT distance="350" swimtime="00:02:28.21" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="28685" number="1" reactiontime="+81" />
                    <RELAYPOSITION athleteid="28696" number="2" reactiontime="+41" />
                    <RELAYPOSITION athleteid="28690" number="3" reactiontime="+59" />
                    <RELAYPOSITION athleteid="27813" number="4" reactiontime="+22" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="15" agetotalmin="14" gender="M" name="Team Saxony HC" number="1">
              <RESULTS>
                <RESULT eventid="26768" reactiontime="+92" swimtime="00:01:37.80" resultid="29390" entrytime="00:01:37.55">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:24.09" />
                    <SPLIT distance="100" swimtime="00:00:50.51" />
                    <SPLIT distance="150" swimtime="00:01:15.81" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="28720" number="1" reactiontime="+92" />
                    <RELAYPOSITION athleteid="28760" number="2" reactiontime="+49" />
                    <RELAYPOSITION athleteid="29213" number="3" reactiontime="+52" />
                    <RELAYPOSITION athleteid="29212" number="4" reactiontime="+95" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="17" agemin="16" agetotalmax="-1" agetotalmin="-1" gender="F" name="Germany DB">
              <RESULTS>
                <RESULT comment="A2 - Niet gestart" eventid="1140" status="DSQ" swimtime="00:00:00.00" resultid="29491" late="yes">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="28721" number="1" status="DSQ" />
                    <RELAYPOSITION athleteid="28702" number="2" status="DSQ" />
                    <RELAYPOSITION athleteid="28722" number="3" status="DSQ" />
                    <RELAYPOSITION athleteid="28707" number="4" status="DSQ" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="15" agetotalmin="14" gender="F" name="Team Saxony DC">
              <RESULTS>
                <RESULT eventid="1217" reactiontime="+97" swimtime="00:03:28.55" resultid="29494" late="yes">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.10" />
                    <SPLIT distance="100" swimtime="00:00:58.31" />
                    <SPLIT distance="150" swimtime="00:01:23.65" />
                    <SPLIT distance="200" swimtime="00:01:51.01" />
                    <SPLIT distance="250" swimtime="00:02:16.85" />
                    <SPLIT distance="300" swimtime="00:02:45.39" />
                    <SPLIT distance="350" swimtime="00:03:05.74" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="28721" number="1" reactiontime="+97" />
                    <RELAYPOSITION athleteid="28702" number="2" reactiontime="+93" />
                    <RELAYPOSITION athleteid="28722" number="3" reactiontime="+60" />
                    <RELAYPOSITION athleteid="28707" number="4" reactiontime="+18" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="15" agetotalmin="14" gender="F" name="Team Saxony2 DC">
              <RESULTS>
                <RESULT eventid="26758" reactiontime="+100" swimtime="00:01:30.97" resultid="29486" late="yes">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:24.37" />
                    <SPLIT distance="100" swimtime="00:00:42.63" />
                    <SPLIT distance="150" swimtime="00:01:08.90" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="28722" number="1" reactiontime="+100" />
                    <RELAYPOSITION athleteid="28707" number="2" />
                    <RELAYPOSITION athleteid="28721" number="3" reactiontime="+89" />
                    <RELAYPOSITION athleteid="28702" number="4" reactiontime="+61" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="15" agetotalmin="14" gender="F" name="Team Saxony 2 DC" number="1">
              <RESULTS>
                <RESULT eventid="1217" reactiontime="+107" swimtime="00:03:17.05" resultid="29395" entrytime="00:03:13.04">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:22.81" />
                    <SPLIT distance="100" swimtime="00:00:47.89" />
                    <SPLIT distance="150" swimtime="00:01:13.48" />
                    <SPLIT distance="200" swimtime="00:01:40.94" />
                    <SPLIT distance="250" swimtime="00:02:04.56" />
                    <SPLIT distance="300" swimtime="00:02:30.60" />
                    <SPLIT distance="350" swimtime="00:02:52.36" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="29263" number="1" reactiontime="+107" />
                    <RELAYPOSITION athleteid="29268" number="2" reactiontime="+89" />
                    <RELAYPOSITION athleteid="28723" number="3" reactiontime="+75" />
                    <RELAYPOSITION athleteid="28713" number="4" reactiontime="+29" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="15" agetotalmin="14" gender="F" name="Team Saxony DC" number="1">
              <RESULTS>
                <RESULT eventid="26758" reactiontime="+106" swimtime="00:01:26.49" resultid="29388" entrytime="00:01:27.23">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:21.70" />
                    <SPLIT distance="100" swimtime="00:00:44.08" />
                    <SPLIT distance="150" swimtime="00:01:06.16" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="29263" number="1" reactiontime="+106" />
                    <RELAYPOSITION athleteid="29268" number="2" reactiontime="+89" />
                    <RELAYPOSITION athleteid="28723" number="3" reactiontime="+71" />
                    <RELAYPOSITION athleteid="28713" number="4" reactiontime="+36" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="34" agetotalmin="18" gender="X" name="Team Saxony GA" number="1">
              <RESULTS>
                <RESULT eventid="1210" reactiontime="+81" swimtime="00:01:11.91" resultid="29393" entrytime="00:01:11.25">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:16.27" />
                    <SPLIT distance="100" swimtime="00:00:35.28" />
                    <SPLIT distance="150" swimtime="00:00:54.38" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="27813" number="1" reactiontime="+81" />
                    <RELAYPOSITION athleteid="28713" number="2" />
                    <RELAYPOSITION athleteid="29263" number="3" />
                    <RELAYPOSITION athleteid="28690" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="17" agemin="16" agetotalmax="-1" agetotalmin="-1" gender="X" name="Team Saxony GB" number="1">
              <RESULTS>
                <RESULT eventid="1140" reactiontime="+85" swimtime="00:03:57.45" resultid="29392" entrytime="00:03:40.06">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.11" />
                    <SPLIT distance="100" swimtime="00:00:57.38" />
                    <SPLIT distance="150" swimtime="00:01:30.81" />
                    <SPLIT distance="200" swimtime="00:02:05.92" />
                    <SPLIT distance="250" swimtime="00:02:35.22" />
                    <SPLIT distance="300" swimtime="00:03:08.89" />
                    <SPLIT distance="350" swimtime="00:03:31.73" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="28696" number="1" reactiontime="+85" />
                    <RELAYPOSITION athleteid="28721" number="2" reactiontime="+101" />
                    <RELAYPOSITION athleteid="28722" number="3" reactiontime="+76" />
                    <RELAYPOSITION athleteid="28690" number="4" reactiontime="+26" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="17" agetotalmin="16" gender="X" name="Team Saxony GB" number="1">
              <RESULTS>
                <RESULT eventid="1210" reactiontime="+99" swimtime="00:01:24.08" resultid="29394" entrytime="00:01:23.52">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:20.63" />
                    <SPLIT distance="100" swimtime="00:00:43.82" />
                    <SPLIT distance="150" swimtime="00:01:05.21" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="28723" number="1" reactiontime="+99" />
                    <RELAYPOSITION athleteid="28720" number="2" reactiontime="+16" />
                    <RELAYPOSITION athleteid="27878" number="3" reactiontime="+66" />
                    <RELAYPOSITION athleteid="28696" number="4" reactiontime="+19" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="15" agemin="14" agetotalmax="-1" agetotalmin="-1" gender="X" name="Team Saxony GC" number="1">
              <RESULTS>
                <RESULT eventid="1140" reactiontime="+78" swimtime="00:03:33.35" resultid="29391" entrytime="00:03:15.73">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:23.66" />
                    <SPLIT distance="100" swimtime="00:00:49.87" />
                    <SPLIT distance="150" swimtime="00:01:17.91" />
                    <SPLIT distance="200" swimtime="00:01:47.29" />
                    <SPLIT distance="250" swimtime="00:02:13.48" />
                    <SPLIT distance="300" swimtime="00:02:43.77" />
                    <SPLIT distance="350" swimtime="00:03:06.96" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="27813" number="1" reactiontime="+78" />
                    <RELAYPOSITION athleteid="28723" number="2" reactiontime="+58" />
                    <RELAYPOSITION athleteid="28713" number="3" reactiontime="+35" />
                    <RELAYPOSITION athleteid="28685" number="4" reactiontime="+15" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="RIESA/DRES" clubid="22879" name="RIESA/DRESDEN" />
        <CLUB type="CLUB" nation="NED" clubid="18186" name="Unattached">
          <COACHES>
            <COACH firstname="Simone" gender="M" lastname="Esch" nameprefix="van" type="HEADCOACH" />
          </COACHES>
          <OFFICIALS>
            <OFFICIAL officialid="21315" firstname="Sven" gender="M" grade="Lijnrechter" lastname="Harteveld" nation="NED" />
            <OFFICIAL officialid="23288" firstname="Simone" gender="F" grade="Ploegleider" lastname="Esch" nameprefix="van" nation="NED" />
            <OFFICIAL officialid="25542" firstname="Mireille" gender="F" grade="Tijdwaarnemer" lastname="Harteveld" nation="NED" />
            <OFFICIAL officialid="21335" firstname="Mireille" gender="F" grade="Speaker" lastname="Harteveld" nation="NED" />
          </OFFICIALS>
        </CLUB>
        <CLUB type="CLUB" code="GAST" nation="NED" clubid="28021" name="Gastzwemmers" shortname="Gast">
          <ATHLETES>
            <ATHLETE firstname="Emese" lastname="Olson" birthdate="2001-05-09" gender="F" nation="NED" license="9265736" athleteid="28105">
              <RESULTS>
                <RESULT comment="A3 - De aangegeven zwemwijze niet uitgevoerd (oa duiken)" eventid="1053" reactiontime="+98" status="DSQ" swimtime="00:00:24.42" resultid="28106" />
                <RESULT eventid="1120" points="501" reactiontime="+85" swimtime="00:00:29.37" resultid="28107" />
                <RESULT eventid="1147" points="424" reactiontime="+128" swimtime="00:00:25.08" resultid="28108" />
                <RESULT eventid="1168" points="506" reactiontime="+90" swimtime="00:01:03.74" resultid="28109">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.53" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="TNAP" nation="FRA" clubid="28826" name="Tours Nage avec palmes" shortname="TNAP">
          <ATHLETES>
            <ATHLETE firstname="Olivier" lastname="Milleville" birthdate="1986-01-02" gender="M" nation="FRA" license="A-03-6092549" athleteid="27050">
              <RESULTS>
                <RESULT eventid="1079" points="830" reactiontime="+87" swimtime="00:00:20.29" resultid="28846" entrytime="00:00:19.04" />
                <RESULT eventid="1114" points="2935" reactiontime="+105" swimtime="00:03:22.30" resultid="28847" entrytime="00:03:17.87">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:23.90" />
                    <SPLIT distance="100" swimtime="00:00:49.72" />
                    <SPLIT distance="150" swimtime="00:01:14.89" />
                    <SPLIT distance="200" swimtime="00:01:40.24" />
                    <SPLIT distance="250" swimtime="00:02:06.30" />
                    <SPLIT distance="300" swimtime="00:02:32.23" />
                    <SPLIT distance="350" swimtime="00:02:57.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1153" points="1039" reactiontime="+88" swimtime="00:00:17.89" resultid="28848" entrytime="00:00:17.78" />
                <RESULT eventid="1190" points="1652" reactiontime="+96" swimtime="00:00:40.15" resultid="28849" entrytime="00:00:39.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:19.26" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Benjamin" lastname="Frehel" birthdate="2004-01-01" gender="M" nation="FRA" license="A-15-680624" athleteid="28828">
              <RESULTS>
                <RESULT eventid="1079" points="595" reactiontime="+93" swimtime="00:00:20.15" resultid="28843" entrytime="00:00:19.89" />
                <RESULT eventid="1127" points="811" reactiontime="+85" swimtime="00:00:21.66" resultid="28844" entrytime="00:00:21.69" />
                <RESULT eventid="1153" points="638" reactiontime="+96" swimtime="00:00:18.36" resultid="28845" entrytime="00:00:17.80" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Arthur" lastname="Castel" birthdate="2002-01-01" gender="M" nation="FRA" license="A-08-392250" athleteid="28827">
              <RESULTS>
                <RESULT eventid="1127" points="670" reactiontime="+91" swimtime="00:00:23.08" resultid="28840" entrytime="00:00:22.00" />
                <RESULT eventid="1175" points="681" reactiontime="+89" swimtime="00:00:52.46" resultid="28841" entrytime="00:00:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1190" points="410" reactiontime="+123" swimtime="00:00:49.16" resultid="28842" entrytime="00:00:52.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:23.79" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <OFFICIALS>
            <OFFICIAL officialid="24572" firstname="Olivier" gender="M" grade="Team Captain" lastname="Milleville" nation="FRA" />
          </OFFICIALS>
        </CLUB>
        <CLUB type="CLUB" code="TCD" nation="GER" clubid="28759" name="TC Delitzsch">
          <ATHLETES>
            <ATHLETE firstname="Pepe Milan" lastname="Becker" birthdate="2011-06-20" gender="M" nation="GER" license="154103000196" athleteid="28760">
              <RESULTS>
                <RESULT eventid="1079" points="718" reactiontime="+93" swimtime="00:00:26.31" resultid="28761" entrytime="00:00:26.15" />
                <RESULT eventid="7271" points="696" reactiontime="+91" swimtime="00:02:37.42" resultid="28762" entrytime="00:02:42.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.01" />
                    <SPLIT distance="100" swimtime="00:01:14.52" />
                    <SPLIT distance="150" swimtime="00:01:57.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1175" points="551" reactiontime="+84" swimtime="00:01:08.73" resultid="28763" entrytime="00:01:13.70">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="7295" points="849" reactiontime="+94" swimtime="00:00:57.50" resultid="28764" entrytime="00:00:59.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1190" points="513" reactiontime="+107" swimtime="00:01:06.85" resultid="28765" entrytime="00:01:05.51">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="24862" points="695" reactiontime="+113" swimtime="00:02:16.38" resultid="28766" entrytime="00:02:14.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.14" />
                    <SPLIT distance="100" swimtime="00:01:05.89" />
                    <SPLIT distance="150" swimtime="00:01:43.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1127" points="719" reactiontime="+99" swimtime="00:00:29.81" resultid="28767" entrytime="00:00:30.90" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <OFFICIALS>
            <OFFICIAL officialid="28804" firstname="Sophie" gender="F" grade="Team Captain" lastname="Niemann" nation="GER" />
          </OFFICIALS>
        </CLUB>
        <CLUB type="CLUB" code="SCHW" nation="GER" clubid="22319" name="TSC Schwandorf" />
        <CLUB type="CLUB" code="MVZZ" nation="NED" clubid="16927" name="MonoVinzz">
          <ATHLETES>
            <ATHLETE firstname="Elma" lastname="Corbijn" birthdate="1973-09-17" gender="F" nation="NED" license="42202" athleteid="28434">
              <RESULTS>
                <RESULT comment="Nieuw Nederlands record" eventid="1093" points="3520" reactiontime="+102" swimtime="00:19:43.21" resultid="28435">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.17" />
                    <SPLIT distance="100" swimtime="00:01:09.24" />
                    <SPLIT distance="150" swimtime="00:01:47.66" />
                    <SPLIT distance="200" swimtime="00:02:26.24" />
                    <SPLIT distance="250" swimtime="00:03:05.47" />
                    <SPLIT distance="300" swimtime="00:03:45.06" />
                    <SPLIT distance="350" swimtime="00:04:24.99" />
                    <SPLIT distance="400" swimtime="00:05:04.82" />
                    <SPLIT distance="450" swimtime="00:05:44.28" />
                    <SPLIT distance="500" swimtime="00:06:23.97" />
                    <SPLIT distance="550" swimtime="00:07:03.72" />
                    <SPLIT distance="600" swimtime="00:07:43.23" />
                    <SPLIT distance="650" swimtime="00:08:23.08" />
                    <SPLIT distance="700" swimtime="00:09:03.04" />
                    <SPLIT distance="750" swimtime="00:09:43.02" />
                    <SPLIT distance="800" swimtime="00:10:22.85" />
                    <SPLIT distance="850" swimtime="00:11:03.40" />
                    <SPLIT distance="900" swimtime="00:11:43.48" />
                    <SPLIT distance="950" swimtime="00:12:23.88" />
                    <SPLIT distance="1000" swimtime="00:13:03.99" />
                    <SPLIT distance="1050" swimtime="00:13:44.25" />
                    <SPLIT distance="1100" swimtime="00:14:24.07" />
                    <SPLIT distance="1150" swimtime="00:15:04.12" />
                    <SPLIT distance="1200" swimtime="00:15:44.94" />
                    <SPLIT distance="1250" swimtime="00:16:25.45" />
                    <SPLIT distance="1300" swimtime="00:17:05.81" />
                    <SPLIT distance="1350" swimtime="00:17:46.88" />
                    <SPLIT distance="1400" swimtime="00:18:27.08" />
                    <SPLIT distance="1450" swimtime="00:19:06.49" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Nieuw Nederlands record" eventid="7254" points="13012" reactiontime="+95" swimtime="00:02:33.05" resultid="28436">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.52" />
                    <SPLIT distance="100" swimtime="00:01:12.62" />
                    <SPLIT distance="150" swimtime="00:01:53.92" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Nederlands record" eventid="7278" points="2123" reactiontime="+109" swimtime="00:05:04.04" resultid="28437">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.03" />
                    <SPLIT distance="100" swimtime="00:01:08.38" />
                    <SPLIT distance="150" swimtime="00:01:47.13" />
                    <SPLIT distance="200" swimtime="00:02:27.31" />
                    <SPLIT distance="250" swimtime="00:03:07.15" />
                    <SPLIT distance="300" swimtime="00:03:46.76" />
                    <SPLIT distance="350" swimtime="00:04:27.02" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Nieuw Nederlands record" eventid="1158" points="2863" reactiontime="+102" swimtime="00:10:33.78" resultid="28438">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.43" />
                    <SPLIT distance="100" swimtime="00:01:08.96" />
                    <SPLIT distance="150" swimtime="00:01:48.07" />
                    <SPLIT distance="200" swimtime="00:02:28.71" />
                    <SPLIT distance="250" swimtime="00:03:09.90" />
                    <SPLIT distance="300" swimtime="00:03:51.14" />
                    <SPLIT distance="350" swimtime="00:04:31.99" />
                    <SPLIT distance="400" swimtime="00:05:13.02" />
                    <SPLIT distance="450" swimtime="00:05:53.87" />
                    <SPLIT distance="500" swimtime="00:06:34.71" />
                    <SPLIT distance="550" swimtime="00:07:15.59" />
                    <SPLIT distance="600" swimtime="00:07:56.13" />
                    <SPLIT distance="650" swimtime="00:08:36.93" />
                    <SPLIT distance="700" swimtime="00:09:17.17" />
                    <SPLIT distance="750" swimtime="00:09:56.39" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Nederlands record" eventid="1168" points="1017" reactiontime="+93" swimtime="00:01:06.09" resultid="28439">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="7287" points="830" reactiontime="+88" swimtime="00:01:04.47" resultid="28440">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="24851" points="867" reactiontime="+95" swimtime="00:02:26.04" resultid="28441">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.29" />
                    <SPLIT distance="100" swimtime="00:01:08.73" />
                    <SPLIT distance="150" swimtime="00:01:49.04" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Xafiera" lastname="Hulst" birthdate="2007-09-05" gender="F" nameprefix="van der" nation="NED" license="9250283" athleteid="28442">
              <RESULTS>
                <RESULT eventid="1053" points="587" reactiontime="+87" swimtime="00:00:24.59" resultid="28443" />
                <RESULT eventid="7254" points="720" reactiontime="+93" swimtime="00:02:13.18" resultid="28444">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.31" />
                    <SPLIT distance="100" swimtime="00:01:03.74" />
                    <SPLIT distance="150" swimtime="00:01:38.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="7278" points="568" reactiontime="+97" swimtime="00:04:32.48" resultid="28445">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.58" />
                    <SPLIT distance="100" swimtime="00:01:02.82" />
                    <SPLIT distance="150" swimtime="00:01:36.83" />
                    <SPLIT distance="200" swimtime="00:02:12.40" />
                    <SPLIT distance="250" swimtime="00:02:48.42" />
                    <SPLIT distance="300" swimtime="00:03:24.35" />
                    <SPLIT distance="350" swimtime="00:03:59.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1147" points="559" reactiontime="+102" swimtime="00:00:23.27" resultid="28446" />
                <RESULT eventid="1168" points="671" reactiontime="+97" swimtime="00:01:00.73" resultid="28447">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="7287" points="566" reactiontime="+107" swimtime="00:00:55.90" resultid="28448">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1182" points="461" reactiontime="+109" swimtime="00:00:57.18" resultid="28449">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.20" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <OFFICIALS>
            <OFFICIAL officialid="1529" firstname="Meindert" grade="Kamprechter" lastname="Boon" nation="NED" />
            <OFFICIAL officialid="21306" firstname="Maikel" gender="M" grade="ETW" lastname="Waart" nameprefix="de" nation="NED" />
            <OFFICIAL officialid="23166" firstname="Liesbeth" gender="F" grade="Secretariaat" lastname="Timmer" nation="NED" />
            <OFFICIAL officialid="1536" firstname="Nancy" gender="F" grade="Ploegleider" lastname="Hoek" nation="NED" />
            <OFFICIAL officialid="1528" firstname="Irene" gender="F" grade="Briefloper" lastname="Glas" nation="NED" />
            <OFFICIAL officialid="1532" firstname="Erik" gender="M" grade="Briefloper" lastname="Glas" nation="NED" />
            <OFFICIAL officialid="18241" firstname="Milo" gender="M" grade="Splash" lastname="Grosz" nation="NED" />
            <OFFICIAL officialid="23160" firstname="Nancy" gender="F" grade="Tijdwaarnemer" lastname="Hoek" nation="NED" />
            <OFFICIAL officialid="7616" firstname="Dennis" gender="M" grade="Secretariaat" lastname="Kap" nation="NED" />
          </OFFICIALS>
        </CLUB>
        <CLUB type="CLUB" code="PAN" nation="FRA" clubid="24484" name="Pays d&apos;Aix Natation" />
        <CLUB type="CLUB" code="TC HARZ" nation="GER" clubid="27874" name="TC Harz">
          <ATHLETES>
            <ATHLETE firstname="Fynn" lastname="Härter" birthdate="2008-01-01" gender="M" nation="GER" license="000389" athleteid="29212">
              <RESULTS>
                <RESULT eventid="1079" points="891" reactiontime="+101" swimtime="00:00:21.52" resultid="29224" entrytime="00:00:22.09" />
                <RESULT eventid="1127" points="772" reactiontime="+94" swimtime="00:00:24.93" resultid="29225" entrytime="00:00:24.50" />
                <RESULT eventid="1153" points="844" reactiontime="+114" swimtime="00:00:19.38" resultid="29226" entrytime="00:00:19.93" />
                <RESULT eventid="7295" points="817" reactiontime="+104" swimtime="00:00:48.59" resultid="29227" entrytime="00:00:49.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:23.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="24862" points="857" reactiontime="+106" swimtime="00:01:51.26" resultid="29228" entrytime="00:01:49.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:24.12" />
                    <SPLIT distance="100" swimtime="00:00:53.00" />
                    <SPLIT distance="150" swimtime="00:01:23.28" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Elisabeth" lastname="Risse" birthdate="2007-06-14" gender="F" nation="GER" license="000390" athleteid="27878">
              <RESULTS>
                <RESULT eventid="1093" points="559" reactiontime="+109" swimtime="00:18:17.02" resultid="29219" entrytime="00:17:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.67" />
                    <SPLIT distance="100" swimtime="00:01:02.23" />
                    <SPLIT distance="150" swimtime="00:01:35.98" />
                    <SPLIT distance="200" swimtime="00:02:09.94" />
                    <SPLIT distance="250" swimtime="00:02:43.95" />
                    <SPLIT distance="300" swimtime="00:03:18.33" />
                    <SPLIT distance="350" swimtime="00:03:52.43" />
                    <SPLIT distance="400" swimtime="00:04:28.19" />
                    <SPLIT distance="450" swimtime="00:05:03.53" />
                    <SPLIT distance="500" swimtime="00:05:39.95" />
                    <SPLIT distance="550" swimtime="00:06:15.46" />
                    <SPLIT distance="600" swimtime="00:06:52.00" />
                    <SPLIT distance="650" swimtime="00:07:27.87" />
                    <SPLIT distance="700" swimtime="00:08:04.46" />
                    <SPLIT distance="750" swimtime="00:08:40.70" />
                    <SPLIT distance="800" swimtime="00:09:17.13" />
                    <SPLIT distance="850" swimtime="00:09:52.57" />
                    <SPLIT distance="900" swimtime="00:10:30.04" />
                    <SPLIT distance="950" swimtime="00:11:06.50" />
                    <SPLIT distance="1000" swimtime="00:11:44.90" />
                    <SPLIT distance="1050" swimtime="00:12:21.72" />
                    <SPLIT distance="1100" swimtime="00:12:59.18" />
                    <SPLIT distance="1150" swimtime="00:13:35.63" />
                    <SPLIT distance="1200" swimtime="00:14:13.73" />
                    <SPLIT distance="1250" swimtime="00:14:50.26" />
                    <SPLIT distance="1300" swimtime="00:15:30.21" />
                    <SPLIT distance="1350" swimtime="00:16:10.28" />
                    <SPLIT distance="1400" swimtime="00:16:50.30" />
                    <SPLIT distance="1450" swimtime="00:17:33.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="7278" points="707" reactiontime="+86" swimtime="00:04:13.29" resultid="29220" entrytime="00:04:07.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.52" />
                    <SPLIT distance="100" swimtime="00:00:57.28" />
                    <SPLIT distance="150" swimtime="00:01:28.95" />
                    <SPLIT distance="200" swimtime="00:02:01.12" />
                    <SPLIT distance="250" swimtime="00:02:34.26" />
                    <SPLIT distance="300" swimtime="00:03:07.76" />
                    <SPLIT distance="350" swimtime="00:03:41.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1158" points="642" reactiontime="+93" swimtime="00:09:02.83" resultid="29221" entrytime="00:08:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.76" />
                    <SPLIT distance="100" swimtime="00:01:00.21" />
                    <SPLIT distance="150" swimtime="00:01:33.35" />
                    <SPLIT distance="200" swimtime="00:02:07.09" />
                    <SPLIT distance="250" swimtime="00:02:40.80" />
                    <SPLIT distance="300" swimtime="00:03:15.34" />
                    <SPLIT distance="350" swimtime="00:03:50.39" />
                    <SPLIT distance="400" swimtime="00:04:24.92" />
                    <SPLIT distance="450" swimtime="00:04:59.73" />
                    <SPLIT distance="500" swimtime="00:05:34.21" />
                    <SPLIT distance="550" swimtime="00:06:09.01" />
                    <SPLIT distance="600" swimtime="00:06:45.43" />
                    <SPLIT distance="650" swimtime="00:07:20.90" />
                    <SPLIT distance="700" swimtime="00:07:56.32" />
                    <SPLIT distance="750" swimtime="00:08:29.92" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="A1 - Bewogen of te vroeg weg bij de start (geen tijd noteren)" eventid="7287" reactiontime="+84" status="DSQ" swimtime="00:00:00.00" resultid="29222" entrytime="00:00:49.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:22.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="24851" points="648" reactiontime="+104" swimtime="00:01:59.36" resultid="29223" entrytime="00:01:51.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.79" />
                    <SPLIT distance="100" swimtime="00:00:55.56" />
                    <SPLIT distance="150" swimtime="00:01:27.02" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jan Henrik" lastname="Hass" birthdate="2004-03-30" gender="M" nation="GER" license="000355" athleteid="27877">
              <RESULTS>
                <RESULT eventid="1079" points="675" reactiontime="+110" swimtime="00:00:19.32" resultid="29216" entrytime="00:00:18.87" />
                <RESULT eventid="7271" points="871" reactiontime="+88" swimtime="00:01:54.08" resultid="29217" entrytime="00:01:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.13" />
                    <SPLIT distance="100" swimtime="00:00:55.76" />
                    <SPLIT distance="150" swimtime="00:01:25.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1127" points="688" reactiontime="+83" swimtime="00:00:22.88" resultid="29218" entrytime="00:00:21.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marnie" lastname="Weißenborn" lastname.en="Weißenborn" birthdate="2008-01-01" gender="F" nation="GER" license="000393" athleteid="27879">
              <RESULTS>
                <RESULT eventid="1053" points="940" reactiontime="+106" swimtime="00:00:21.86" resultid="29229" entrytime="00:00:21.60" />
                <RESULT eventid="7254" points="1014" reactiontime="+89" swimtime="00:02:06.14" resultid="29230" entrytime="00:02:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.36" />
                    <SPLIT distance="100" swimtime="00:01:01.04" />
                    <SPLIT distance="150" swimtime="00:01:34.38" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="A2 - Niet gestart" eventid="1120" status="DSQ" swimtime="00:00:00.00" resultid="29231" entrytime="00:00:24.50" />
                <RESULT eventid="1147" points="820" reactiontime="+101" swimtime="00:00:20.52" resultid="29232" entrytime="00:00:19.50" />
                <RESULT eventid="1158" points="782" reactiontime="+112" swimtime="00:08:51.44" resultid="29233" entrytime="00:08:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.05" />
                    <SPLIT distance="100" swimtime="00:01:00.43" />
                    <SPLIT distance="150" swimtime="00:01:33.77" />
                    <SPLIT distance="200" swimtime="00:02:07.45" />
                    <SPLIT distance="250" swimtime="00:02:42.15" />
                    <SPLIT distance="300" swimtime="00:03:15.74" />
                    <SPLIT distance="350" swimtime="00:03:49.97" />
                    <SPLIT distance="400" swimtime="00:04:24.03" />
                    <SPLIT distance="450" swimtime="00:04:58.52" />
                    <SPLIT distance="500" swimtime="00:05:32.82" />
                    <SPLIT distance="550" swimtime="00:06:06.56" />
                    <SPLIT distance="600" swimtime="00:06:40.84" />
                    <SPLIT distance="650" swimtime="00:07:14.32" />
                    <SPLIT distance="700" swimtime="00:07:48.07" />
                    <SPLIT distance="750" swimtime="00:08:21.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="7287" points="986" reactiontime="+107" swimtime="00:00:47.47" resultid="29234" entrytime="00:00:46.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:22.79" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Noah" lastname="Dalichow" birthdate="2003-06-25" gender="M" nation="GER" license="000329" athleteid="27876">
              <RESULTS>
                <RESULT eventid="1079" points="714" reactiontime="+102" swimtime="00:00:18.96" resultid="29214" entrytime="00:00:18.72" />
                <RESULT eventid="1127" points="749" reactiontime="+89" swimtime="00:00:22.24" resultid="29215" entrytime="00:00:21.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Matty" lastname="Schmidt" birthdate="2009-01-01" gender="M" nation="GER" license="000382" athleteid="29213">
              <RESULTS>
                <RESULT eventid="1079" points="547" reactiontime="+101" swimtime="00:00:25.32" resultid="29239" entrytime="00:00:24.87" />
                <RESULT comment="A11 - Uitrusting voldoet niet aan de geldende eisen" eventid="7264" reactiontime="+101" status="DSQ" swimtime="00:00:00.00" resultid="29240" entrytime="00:04:23.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.17" />
                    <SPLIT distance="100" swimtime="00:01:03.92" />
                    <SPLIT distance="150" swimtime="00:01:37.48" />
                    <SPLIT distance="200" swimtime="00:02:12.79" />
                    <SPLIT distance="250" swimtime="00:02:45.17" />
                    <SPLIT distance="300" swimtime="00:03:19.11" />
                    <SPLIT distance="350" swimtime="00:03:52.78" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="C1 - Niet de gehele afstand met het gezicht onder water afgelegd" eventid="1153" reactiontime="+105" status="DSQ" swimtime="00:00:00.00" resultid="29241" entrytime="00:00:26.00" />
                <RESULT eventid="7295" status="WDR" swimtime="00:00:00.00" resultid="29242" entrytime="00:00:55.80" />
                <RESULT eventid="24862" status="WDR" swimtime="00:00:00.00" resultid="29243" entrytime="00:02:00.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marlene" lastname="Zündel" birthdate="2009-09-22" gender="F" nation="GER" license="000391" athleteid="27880">
              <RESULTS>
                <RESULT eventid="7278" points="702" reactiontime="+115" swimtime="00:04:20.44" resultid="29235" entrytime="00:04:19.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.69" />
                    <SPLIT distance="100" swimtime="00:00:59.49" />
                    <SPLIT distance="150" swimtime="00:01:33.08" />
                    <SPLIT distance="200" swimtime="00:02:07.06" />
                    <SPLIT distance="250" swimtime="00:02:39.91" />
                    <SPLIT distance="300" swimtime="00:03:14.01" />
                    <SPLIT distance="350" swimtime="00:03:48.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1158" points="564" reactiontime="+108" swimtime="00:09:52.67" resultid="29236" entrytime="00:09:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.12" />
                    <SPLIT distance="100" swimtime="00:01:04.39" />
                    <SPLIT distance="150" swimtime="00:01:39.96" />
                    <SPLIT distance="200" swimtime="00:02:16.74" />
                    <SPLIT distance="250" swimtime="00:02:51.19" />
                    <SPLIT distance="300" swimtime="00:03:27.92" />
                    <SPLIT distance="350" swimtime="00:04:05.34" />
                    <SPLIT distance="400" swimtime="00:04:41.99" />
                    <SPLIT distance="450" swimtime="00:05:19.86" />
                    <SPLIT distance="500" swimtime="00:05:59.17" />
                    <SPLIT distance="550" swimtime="00:06:39.20" />
                    <SPLIT distance="600" swimtime="00:07:16.99" />
                    <SPLIT distance="650" swimtime="00:07:57.89" />
                    <SPLIT distance="700" swimtime="00:08:37.47" />
                    <SPLIT distance="750" swimtime="00:09:14.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="7287" points="712" reactiontime="+104" swimtime="00:00:52.92" resultid="29237" entrytime="00:00:51.44">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="24851" points="680" reactiontime="+107" swimtime="00:02:00.53" resultid="29238" entrytime="00:01:57.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.86" />
                    <SPLIT distance="100" swimtime="00:00:57.27" />
                    <SPLIT distance="150" swimtime="00:01:29.17" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="34" agetotalmin="18" gender="M" name="TC Harz HA" number="1">
              <RESULTS>
                <RESULT eventid="26768" reactiontime="+97" swimtime="00:01:25.27" resultid="29244" entrytime="00:01:17.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:18.81" />
                    <SPLIT distance="100" swimtime="00:00:37.71" />
                    <SPLIT distance="150" swimtime="00:01:00.03" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="27876" number="1" reactiontime="+97" />
                    <RELAYPOSITION athleteid="27877" number="2" reactiontime="+48" />
                    <RELAYPOSITION athleteid="29212" number="3" reactiontime="+76" />
                    <RELAYPOSITION athleteid="29213" number="4" reactiontime="+87" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="34" agemin="18" agetotalmax="-1" agetotalmin="-1" gender="X">
              <RESULTS>
                <RESULT eventid="1140" reactiontime="+89" swimtime="00:03:34.02" resultid="29489" late="yes">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:23.42" />
                    <SPLIT distance="100" swimtime="00:00:48.75" />
                    <SPLIT distance="150" swimtime="00:01:14.75" />
                    <SPLIT distance="200" swimtime="00:01:43.82" />
                    <SPLIT distance="250" swimtime="00:02:12.06" />
                    <SPLIT distance="300" swimtime="00:02:43.60" />
                    <SPLIT distance="350" swimtime="00:03:07.31" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="27876" number="1" reactiontime="+89" />
                    <RELAYPOSITION athleteid="27879" number="2" reactiontime="+78" />
                    <RELAYPOSITION athleteid="27880" number="3" reactiontime="+34" />
                    <RELAYPOSITION athleteid="27877" number="4" reactiontime="+48" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="34" agemin="18" agetotalmax="-1" agetotalmin="-1" gender="X" name="TC Harz GA" number="1">
              <RESULTS>
                <RESULT comment="A2 - Niet gestart" eventid="1140" status="DSQ" swimtime="00:00:00.00" resultid="29245" entrytime="00:03:40.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="29212" number="1" status="DSQ" />
                    <RELAYPOSITION athleteid="29213" number="2" status="DSQ" />
                    <RELAYPOSITION athleteid="27879" number="3" status="DSQ" />
                    <RELAYPOSITION athleteid="27880" number="4" status="DSQ" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="15" agetotalmin="14" gender="X" name="TC Harz GC" number="1">
              <RESULTS>
                <RESULT comment="C1 - Niet de gehele afstand met het gezicht onder water afgelegd, C1 2e zwemmer, niet gefinisht" eventid="1210" reactiontime="+102" status="DSQ" swimtime="00:00:00.00" resultid="29246" entrytime="00:01:26.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:21.33" />
                    <SPLIT distance="100" swimtime="00:00:48.97" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="27879" number="1" reactiontime="+102" status="DSQ" />
                    <RELAYPOSITION athleteid="29213" number="2" reactiontime="+51" status="DSQ" />
                    <RELAYPOSITION athleteid="27880" number="3" status="DSQ" />
                    <RELAYPOSITION athleteid="29212" number="4" status="DSQ" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
          <OFFICIALS>
            <OFFICIAL officialid="29211" firstname="Holger" gender="M" grade="Team Captain" lastname="Dalichow" nation="GER" />
            <OFFICIAL officialid="27875" firstname="Birgit" gender="F" grade="Team Captain" lastname="Galler" nation="GER" />
          </OFFICIALS>
        </CLUB>
        <CLUB type="CLUB" code="GRASM" nation="BEL" clubid="24777" name="GRASM" />
        <CLUB type="CLUB" code="DRB" nation="NED" clubid="25223" name="Dordtse Reddingsbrigade" shortname="Dordtse RB">
          <OFFICIALS>
            <OFFICIAL officialid="25537" firstname="Sandra" gender="F" grade="Tijdwaarnemer" lastname="Lohuizen" nameprefix="van" nation="NED" />
          </OFFICIALS>
        </CLUB>
        <CLUB type="CLUB" code="TC NAUTILU" nation="GER" clubid="26032" name="TC Nautilus Mitterteich" shortname="TC Nautilus">
          <OFFICIALS>
            <OFFICIAL officialid="26642" firstname="Roman" gender="M" grade="Team Captain" lastname="Heinrich" nation="GER" />
          </OFFICIALS>
        </CLUB>
        <CLUB type="CLUB" code="TSCW" nation="GER" clubid="26996" name="TSC Weimar">
          <OFFICIALS>
            <OFFICIAL officialid="27685" firstname="Monique" gender="F" grade="Team Captain" lastname="Klabunde - de Jager" nation="GER" />
          </OFFICIALS>
        </CLUB>
        <CLUB type="CLUB" code="PFNAP" nation="FRA" clubid="27806" name="PF NAP AIX" shortname="PFNAP">
          <ATHLETES>
            <ATHLETE firstname="Maïwenn" lastname="Hamon" birthdate="2003-08-11" gender="F" nation="FRA" license="A-15-691710" athleteid="27808">
              <RESULTS>
                <RESULT comment="A3 - De aangegeven zwemwijze niet uitgevoerd (oa duiken)" eventid="1053" reactiontime="+92" status="DSQ" swimtime="00:00:18.94" resultid="28792" entrytime="00:00:18.30" />
                <RESULT eventid="1120" points="934" reactiontime="+79" swimtime="00:00:23.86" resultid="28793" entrytime="00:00:23.50" />
                <RESULT comment="Backup tijd" eventid="1147" points="1271" reactiontime="+89" swimtime="00:00:17.40" resultid="28794" entrytime="00:00:16.99" />
                <RESULT eventid="7287" status="WDR" swimtime="00:00:00.00" resultid="28795" entrytime="00:00:38.10" />
                <RESULT eventid="1182" points="1123" reactiontime="+100" swimtime="00:00:42.50" resultid="29485">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:19.64" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Colas" lastname="Zugmeyer" birthdate="2001-03-11" gender="M" nation="FRA" license="A-12-557961" athleteid="28784">
              <RESULTS>
                <RESULT eventid="1079" points="1068" reactiontime="+86" swimtime="00:00:16.58" resultid="28787" entrytime="00:00:15.87" />
                <RESULT eventid="7264" points="1059" reactiontime="+92" swimtime="00:03:12.73" resultid="28788" entrytime="00:03:05.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:22.58" />
                    <SPLIT distance="100" swimtime="00:00:46.77" />
                    <SPLIT distance="150" swimtime="00:01:11.24" />
                    <SPLIT distance="200" swimtime="00:01:35.94" />
                    <SPLIT distance="250" swimtime="00:02:00.61" />
                    <SPLIT distance="300" swimtime="00:02:25.62" />
                    <SPLIT distance="350" swimtime="00:02:49.50" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Backup tijd" eventid="1153" points="946" reactiontime="+84" swimtime="00:00:16.10" resultid="28789" entrytime="00:00:15.49" />
                <RESULT eventid="7295" points="1176" reactiontime="+86" swimtime="00:00:37.34" resultid="28790" entrytime="00:00:36.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:18.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1190" points="989" reactiontime="+100" swimtime="00:00:36.67" resultid="28791" entrytime="00:00:35.01">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:17.77" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Adrien" lastname="Ghirardi" birthdate="1997-07-12" gender="M" nation="FRA" license="A-18-797886" athleteid="28786">
              <RESULTS>
                <RESULT eventid="7271" points="1079" reactiontime="+79" swimtime="00:01:46.24" resultid="28800" entrytime="00:01:40.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:24.53" />
                    <SPLIT distance="100" swimtime="00:00:52.21" />
                    <SPLIT distance="150" swimtime="00:01:20.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1127" points="983" reactiontime="+77" swimtime="00:00:20.31" resultid="28801" entrytime="00:00:19.92" />
                <RESULT eventid="1175" points="1125" reactiontime="+80" swimtime="00:00:44.37" resultid="28802" entrytime="00:00:43.16">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:20.74" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ewen" lastname="Hamon" birthdate="2005-08-01" gender="M" nation="FRA" license="A-16-742345" athleteid="28785">
              <RESULTS>
                <RESULT eventid="1079" points="1028" reactiontime="+81" swimtime="00:00:16.79" resultid="28796" entrytime="00:00:17.10" />
                <RESULT comment="A1 - Bewogen of te vroeg weg bij de start (geen tijd noteren)" eventid="1153" reactiontime="+51" status="DSQ" swimtime="00:00:00.00" resultid="28797" entrytime="00:00:15.97" />
                <RESULT eventid="1190" points="928" reactiontime="+100" swimtime="00:00:37.46" resultid="28798" entrytime="00:00:35.40">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:18.51" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <OFFICIALS>
            <OFFICIAL officialid="27807" firstname="Cyril" gender="M" grade="Team Captain" lastname="Aoubid" nation="FRA" />
          </OFFICIALS>
        </CLUB>
        <CLUB type="CLUB" code="TCSP" nation="GER" clubid="26139" name="TC Submarin Pössneck" shortname="TCSP">
          <COACHES>
            <COACH firstname="Daniela" gender="F" lastname="Matthes" nation="GER" type="COACH" />
          </COACHES>
          <OFFICIALS>
            <OFFICIAL officialid="26155" firstname="Daniela" gender="F" grade="Team Captain" lastname="Matthes" nation="GER" />
          </OFFICIALS>
        </CLUB>
        <CLUB type="CLUB" code="DUC" nation="GER" clubid="23168" name="DUC Darmstadt" shortname="DUC">
          <OFFICIALS>
            <OFFICIAL officialid="23169" firstname="Frank" gender="M" grade="Tijdwaarnemer" lastname="Spieß" nation="GER" license="DLD 50" />
            <OFFICIAL officialid="23167" firstname="Tassilo" gender="M" grade="Tijdwaarnemer" lastname="Arndt" nation="GER" license="DLD 654" />
          </OFFICIALS>
        </CLUB>
        <CLUB type="CLUB" code="CSAKB" nation="FRA" clubid="26021" name="CSA Kremlin-Bicetre" shortname="CSA KB">
          <ATHLETES>
            <ATHLETE firstname="Clara" lastname="Real" birthdate="2004-01-01" gender="F" nation="FRA" license="A-19-834976" athleteid="28825">
              <RESULTS>
                <RESULT eventid="1053" points="804" reactiontime="+100" swimtime="00:00:21.46" resultid="28833" entrytime="00:00:20.88" />
                <RESULT eventid="1147" points="950" reactiontime="+96" swimtime="00:00:19.17" resultid="28834" entrytime="00:00:18.61" />
                <RESULT eventid="1182" points="1008" reactiontime="+106" swimtime="00:00:44.06" resultid="28835" entrytime="00:00:42.89">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:21.36" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Evan" lastname="Morin" birthdate="2006-07-22" gender="M" nation="FRA" license="A-16-720818" athleteid="27055">
              <RESULTS>
                <RESULT eventid="7271" points="1303" reactiontime="+96" swimtime="00:01:42.96" resultid="28836" entrytime="00:01:48.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:23.82" />
                    <SPLIT distance="100" swimtime="00:00:49.86" />
                    <SPLIT distance="150" swimtime="00:01:16.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1127" points="1112" reactiontime="+92" swimtime="00:00:21.82" resultid="28837" entrytime="00:00:22.00" />
                <RESULT eventid="1175" points="1193" reactiontime="+88" swimtime="00:00:47.32" resultid="28838" entrytime="00:00:48.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:23.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1203" points="1261" reactiontime="+99" swimtime="00:03:40.03" resultid="28839" entrytime="00:03:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:24.46" />
                    <SPLIT distance="100" swimtime="00:00:51.28" />
                    <SPLIT distance="150" swimtime="00:01:19.40" />
                    <SPLIT distance="200" swimtime="00:01:47.79" />
                    <SPLIT distance="250" swimtime="00:02:16.07" />
                    <SPLIT distance="300" swimtime="00:02:44.79" />
                    <SPLIT distance="350" swimtime="00:03:13.32" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <OFFICIALS>
            <OFFICIAL officialid="26640" firstname="Valérie" gender="F" grade="Team Captain" lastname="Morin" nation="FRA" />
            <OFFICIAL officialid="28824" firstname="Olivier" gender="M" grade="Team Captain" lastname="Milleville" nation="FRA" />
            <OFFICIAL officialid="27684" firstname="Alex" gender="M" grade="Team Captain" lastname="Neumann" nation="FRA" />
          </OFFICIALS>
        </CLUB>
        <CLUB type="CLUB" code="HSTSG" nation="GER" clubid="26170" name="Hochschul Tauchsportgruppe" shortname="HSTSG" />
        <CLUB type="CLUB" code="TCH" nation="GER" clubid="22014" name="Tauchclub Heilbronn">
          <ATHLETES>
            <ATHLETE firstname="Leona" lastname="Ruedel" birthdate="2004-07-28" gender="F" nation="GER" license="124012000739" athleteid="27536">
              <RESULTS>
                <RESULT eventid="1053" points="778" reactiontime="+91" swimtime="00:00:21.70" resultid="28520" entrytime="00:00:21.52" />
                <RESULT eventid="7278" points="853" reactiontime="+101" swimtime="00:03:56.31" resultid="28521" entrytime="00:03:55.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.71" />
                    <SPLIT distance="100" swimtime="00:00:54.10" />
                    <SPLIT distance="150" swimtime="00:01:24.42" />
                    <SPLIT distance="200" swimtime="00:01:55.44" />
                    <SPLIT distance="250" swimtime="00:02:26.74" />
                    <SPLIT distance="300" swimtime="00:02:57.73" />
                    <SPLIT distance="350" swimtime="00:03:28.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1147" points="848" reactiontime="+98" swimtime="00:00:19.91" resultid="28522" entrytime="00:00:19.14" />
                <RESULT eventid="7287" points="882" reactiontime="+91" swimtime="00:00:47.87" resultid="28523" entrytime="00:00:46.67">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:23.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1182" points="760" reactiontime="+110" swimtime="00:00:48.41" resultid="28524" entrytime="00:00:45.83">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:23.80" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Benedikt" lastname="Bilicz" birthdate="2007-08-28" gender="M" nation="GER" license="124012000783" athleteid="27505">
              <RESULTS>
                <RESULT eventid="1079" points="870" reactiontime="+97" swimtime="00:00:19.63" resultid="28530" entrytime="00:00:19.76" />
                <RESULT eventid="7264" points="698" reactiontime="+97" swimtime="00:03:56.70" resultid="28531" entrytime="00:03:54.18">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:23.45" />
                    <SPLIT distance="100" swimtime="00:00:50.85" />
                    <SPLIT distance="150" swimtime="00:01:19.97" />
                    <SPLIT distance="200" swimtime="00:01:51.47" />
                    <SPLIT distance="250" swimtime="00:02:23.89" />
                    <SPLIT distance="300" swimtime="00:02:56.28" />
                    <SPLIT distance="350" swimtime="00:03:28.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1153" points="998" reactiontime="+96" swimtime="00:00:16.96" resultid="28532" entrytime="00:00:17.22" />
                <RESULT eventid="7295" points="819" reactiontime="+93" swimtime="00:00:43.63" resultid="28533" entrytime="00:00:45.07">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:20.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="24862" points="850" reactiontime="+93" swimtime="00:01:48.25" resultid="28534" entrytime="00:01:45.07">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:23.44" />
                    <SPLIT distance="100" swimtime="00:00:50.59" />
                    <SPLIT distance="150" swimtime="00:01:19.47" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Hannah" lastname="Grimm" birthdate="2008-04-18" gender="F" nation="GER" license="1204012000800" athleteid="27512">
              <RESULTS>
                <RESULT eventid="1053" points="703" reactiontime="+109" swimtime="00:00:24.08" resultid="28504" entrytime="00:00:23.81" />
                <RESULT eventid="7278" points="549" reactiontime="+106" swimtime="00:04:42.66" resultid="28505" entrytime="00:04:41.88">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.69" />
                    <SPLIT distance="100" swimtime="00:01:04.86" />
                    <SPLIT distance="150" swimtime="00:01:41.34" />
                    <SPLIT distance="200" swimtime="00:02:18.25" />
                    <SPLIT distance="250" swimtime="00:02:55.51" />
                    <SPLIT distance="300" swimtime="00:03:33.10" />
                    <SPLIT distance="350" swimtime="00:04:09.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1147" points="631" reactiontime="+123" swimtime="00:00:22.39" resultid="28506" entrytime="00:00:22.58" />
                <RESULT eventid="7287" points="676" reactiontime="+108" swimtime="00:00:53.84" resultid="28507" entrytime="00:00:54.32">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="24851" points="573" reactiontime="+122" swimtime="00:02:07.60" resultid="28508" entrytime="00:02:07.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.16" />
                    <SPLIT distance="100" swimtime="00:01:01.77" />
                    <SPLIT distance="150" swimtime="00:01:35.23" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Tobias" lastname="Fabriz" birthdate="2003-06-19" gender="M" nation="GER" license="124012000686" athleteid="27507">
              <RESULTS>
                <RESULT eventid="1079" points="695" reactiontime="+105" swimtime="00:00:19.13" resultid="28535" entrytime="00:00:19.21" />
                <RESULT eventid="1153" points="842" reactiontime="+95" swimtime="00:00:16.74" resultid="28536" entrytime="00:00:17.05" />
                <RESULT eventid="7295" points="729" reactiontime="+95" swimtime="00:00:43.78" resultid="28537" entrytime="00:00:42.93">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:20.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1190" points="648" reactiontime="+108" swimtime="00:00:42.21" resultid="28538" entrytime="00:00:41.65">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:20.29" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Beeke Alea" lastname="Phillipp" birthdate="2004-12-28" gender="F" nation="GER" license="124012000694" athleteid="27524">
              <RESULTS>
                <RESULT eventid="1053" points="803" reactiontime="+116" swimtime="00:00:21.47" resultid="28515" entrytime="00:00:21.23" />
                <RESULT eventid="7278" points="855" reactiontime="+99" swimtime="00:03:56.07" resultid="28516" entrytime="00:03:58.38">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:24.95" />
                    <SPLIT distance="100" swimtime="00:00:52.42" />
                    <SPLIT distance="150" swimtime="00:01:21.65" />
                    <SPLIT distance="200" swimtime="00:01:51.90" />
                    <SPLIT distance="250" swimtime="00:02:22.59" />
                    <SPLIT distance="300" swimtime="00:02:53.78" />
                    <SPLIT distance="350" swimtime="00:03:25.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1147" points="853" reactiontime="+98" swimtime="00:00:19.87" resultid="28517" entrytime="00:00:19.27" />
                <RESULT eventid="7287" points="876" reactiontime="+96" swimtime="00:00:47.98" resultid="28518" entrytime="00:00:46.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:22.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1182" points="871" reactiontime="+118" swimtime="00:00:46.26" resultid="28519" entrytime="00:00:45.53">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:22.11" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Frida" lastname="Leleux" birthdate="2012-01-01" gender="F" nation="GER" license="124012000862" athleteid="28488">
              <RESULTS>
                <RESULT eventid="1053" points="836" reactiontime="+129" swimtime="00:00:27.26" resultid="28489" entrytime="00:00:26.01" />
                <RESULT eventid="7278" points="837" reactiontime="+128" swimtime="00:05:25.51" resultid="28490" entrytime="00:05:11.34">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.84" />
                    <SPLIT distance="100" swimtime="00:01:14.75" />
                    <SPLIT distance="150" swimtime="00:01:58.02" />
                    <SPLIT distance="200" swimtime="00:02:40.90" />
                    <SPLIT distance="250" swimtime="00:03:23.41" />
                    <SPLIT distance="300" swimtime="00:04:08.38" />
                    <SPLIT distance="350" swimtime="00:04:50.39" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Backup tijd" eventid="1168" points="711" reactiontime="+107" swimtime="00:01:12.27" resultid="28491" entrytime="00:01:02.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="7287" points="942" reactiontime="+103" swimtime="00:01:00.16" resultid="28492" entrytime="00:01:00.68">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="24851" points="832" reactiontime="+119" swimtime="00:02:20.50" resultid="28493" entrytime="00:02:18.33">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.39" />
                    <SPLIT distance="100" swimtime="00:01:09.46" />
                    <SPLIT distance="150" swimtime="00:01:47.93" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Sina" lastname="Rettig" birthdate="2009-02-07" gender="F" nation="GER" license="124012000773" athleteid="27530">
              <RESULTS>
                <RESULT eventid="1053" points="631" reactiontime="+105" swimtime="00:00:24.97" resultid="28494" entrytime="00:00:24.69" />
                <RESULT eventid="7278" points="541" reactiontime="+98" swimtime="00:04:43.98" resultid="28495" entrytime="00:05:00.78">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.82" />
                    <SPLIT distance="100" swimtime="00:01:04.34" />
                    <SPLIT distance="150" swimtime="00:01:40.58" />
                    <SPLIT distance="200" swimtime="00:02:19.30" />
                    <SPLIT distance="250" swimtime="00:02:57.34" />
                    <SPLIT distance="300" swimtime="00:03:34.93" />
                    <SPLIT distance="350" swimtime="00:04:10.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1147" points="451" reactiontime="+116" swimtime="00:00:25.04" resultid="28496" entrytime="00:00:23.77" />
                <RESULT eventid="7287" points="614" reactiontime="+103" swimtime="00:00:55.60" resultid="28497" entrytime="00:00:56.78">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="24851" points="482" reactiontime="+109" swimtime="00:02:15.20" resultid="28498" entrytime="00:02:10.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.50" />
                    <SPLIT distance="100" swimtime="00:01:05.53" />
                    <SPLIT distance="150" swimtime="00:01:42.14" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Esther-Sophie" lastname="Seidel" birthdate="2008-11-07" gender="F" nation="GER" license="124012000774" athleteid="27542">
              <RESULTS>
                <RESULT eventid="1053" points="857" reactiontime="+123" swimtime="00:00:22.55" resultid="28509" entrytime="00:00:21.92" />
                <RESULT eventid="7278" points="682" reactiontime="+122" swimtime="00:04:22.90" resultid="28510" entrytime="00:04:26.11">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.13" />
                    <SPLIT distance="100" swimtime="00:01:02.20" />
                    <SPLIT distance="150" swimtime="00:01:36.17" />
                    <SPLIT distance="200" swimtime="00:02:10.56" />
                    <SPLIT distance="250" swimtime="00:02:44.93" />
                    <SPLIT distance="300" swimtime="00:03:19.45" />
                    <SPLIT distance="350" swimtime="00:03:53.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1147" points="725" reactiontime="+114" swimtime="00:00:21.38" resultid="28511" entrytime="00:00:20.77" />
                <RESULT eventid="1158" points="657" reactiontime="+114" swimtime="00:09:23.13" resultid="28512" entrytime="00:09:43.45">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.22" />
                    <SPLIT distance="100" swimtime="00:01:02.71" />
                    <SPLIT distance="150" swimtime="00:01:37.82" />
                    <SPLIT distance="200" swimtime="00:02:14.48" />
                    <SPLIT distance="250" swimtime="00:02:50.35" />
                    <SPLIT distance="300" swimtime="00:03:28.08" />
                    <SPLIT distance="350" swimtime="00:04:04.78" />
                    <SPLIT distance="400" swimtime="00:04:42.40" />
                    <SPLIT distance="450" swimtime="00:05:18.32" />
                    <SPLIT distance="500" swimtime="00:05:55.33" />
                    <SPLIT distance="550" swimtime="00:06:32.68" />
                    <SPLIT distance="600" swimtime="00:07:10.03" />
                    <SPLIT distance="650" swimtime="00:07:47.60" />
                    <SPLIT distance="700" swimtime="00:08:22.78" />
                    <SPLIT distance="750" swimtime="00:08:54.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="24851" points="680" reactiontime="+118" swimtime="00:02:00.53" resultid="28514" entrytime="00:01:58.57">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.34" />
                    <SPLIT distance="100" swimtime="00:00:57.34" />
                    <SPLIT distance="150" swimtime="00:01:30.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="7287" points="792" reactiontime="+112" swimtime="00:00:51.07" resultid="28769" entrytime="00:00:50.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:24.30" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Elisa" lastname="Hölzer" birthdate="2009-10-19" gender="F" nation="GER" license="124012000775" athleteid="27506">
              <RESULTS>
                <RESULT eventid="1053" points="767" reactiontime="+99" swimtime="00:00:23.40" resultid="28499" entrytime="00:00:23.27" />
                <RESULT eventid="7278" points="740" reactiontime="+105" swimtime="00:04:15.86" resultid="28500" entrytime="00:04:17.15">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.21" />
                    <SPLIT distance="100" swimtime="00:00:57.58" />
                    <SPLIT distance="150" swimtime="00:01:30.49" />
                    <SPLIT distance="200" swimtime="00:02:04.44" />
                    <SPLIT distance="250" swimtime="00:02:38.49" />
                    <SPLIT distance="300" swimtime="00:03:12.29" />
                    <SPLIT distance="350" swimtime="00:03:44.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1147" points="652" reactiontime="+103" swimtime="00:00:22.15" resultid="28501" entrytime="00:00:22.08" />
                <RESULT eventid="7287" points="808" reactiontime="+102" swimtime="00:00:50.73" resultid="28502" entrytime="00:00:51.34">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:24.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="24851" points="728" reactiontime="+104" swimtime="00:01:57.80" resultid="28503" entrytime="00:01:56.18">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.99" />
                    <SPLIT distance="100" swimtime="00:00:56.30" />
                    <SPLIT distance="150" swimtime="00:01:27.85" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Elias" lastname="Korb" birthdate="2011-02-28" gender="M" nation="GER" license="124012000790" athleteid="27518">
              <RESULTS>
                <RESULT eventid="1079" points="839" reactiontime="+117" swimtime="00:00:24.99" resultid="28525" entrytime="00:00:25.89" />
                <RESULT eventid="7264" points="1280" reactiontime="+118" swimtime="00:04:10.07" resultid="28526" entrytime="00:04:14.93">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.94" />
                    <SPLIT distance="100" swimtime="00:00:59.19" />
                    <SPLIT distance="150" swimtime="00:01:31.70" />
                    <SPLIT distance="200" swimtime="00:02:04.25" />
                    <SPLIT distance="250" swimtime="00:02:37.35" />
                    <SPLIT distance="300" swimtime="00:03:10.68" />
                    <SPLIT distance="350" swimtime="00:03:42.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="16574" points="1115" reactiontime="+129" swimtime="00:08:51.06" resultid="28527" entrytime="00:10:37.32">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.38" />
                    <SPLIT distance="100" swimtime="00:01:02.33" />
                    <SPLIT distance="150" swimtime="00:01:35.96" />
                    <SPLIT distance="200" swimtime="00:02:09.64" />
                    <SPLIT distance="250" swimtime="00:02:44.13" />
                    <SPLIT distance="300" swimtime="00:03:19.20" />
                    <SPLIT distance="350" swimtime="00:03:52.91" />
                    <SPLIT distance="400" swimtime="00:04:26.71" />
                    <SPLIT distance="450" swimtime="00:05:00.70" />
                    <SPLIT distance="500" swimtime="00:05:34.96" />
                    <SPLIT distance="550" swimtime="00:06:09.03" />
                    <SPLIT distance="600" swimtime="00:06:42.61" />
                    <SPLIT distance="650" swimtime="00:07:16.36" />
                    <SPLIT distance="700" swimtime="00:07:50.12" />
                    <SPLIT distance="750" swimtime="00:08:22.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="7295" points="896" reactiontime="+120" swimtime="00:00:56.49" resultid="28528" entrytime="00:00:56.77">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="24862" points="866" reactiontime="+114" swimtime="00:02:06.76" resultid="28529" entrytime="00:02:01.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.78" />
                    <SPLIT distance="100" swimtime="00:01:01.78" />
                    <SPLIT distance="150" swimtime="00:01:36.14" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="15" agetotalmin="14" gender="F" name="TC Heilbronn 2 DC" number="1">
              <RESULTS>
                <RESULT eventid="26758" reactiontime="+103" swimtime="00:01:34.25" resultid="28540" entrytime="00:01:34.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:23.53" />
                    <SPLIT distance="100" swimtime="00:00:48.94" />
                    <SPLIT distance="150" swimtime="00:01:12.65" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="27512" number="1" reactiontime="+103" />
                    <RELAYPOSITION athleteid="27530" number="2" reactiontime="+87" />
                    <RELAYPOSITION athleteid="27506" number="3" reactiontime="+79" />
                    <RELAYPOSITION athleteid="27542" number="4" reactiontime="+87" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="15" agetotalmin="14" gender="F" name="TC Heilbronn 3 DC" number="1">
              <RESULTS>
                <RESULT eventid="1217" reactiontime="+110" swimtime="00:03:41.10" resultid="28541" entrytime="00:03:34.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.10" />
                    <SPLIT distance="100" swimtime="00:00:53.47" />
                    <SPLIT distance="150" swimtime="00:01:21.35" />
                    <SPLIT distance="200" swimtime="00:01:53.81" />
                    <SPLIT distance="250" swimtime="00:02:21.12" />
                    <SPLIT distance="300" swimtime="00:02:50.27" />
                    <SPLIT distance="350" swimtime="00:03:13.93" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="27506" number="1" reactiontime="+110" />
                    <RELAYPOSITION athleteid="27530" number="2" reactiontime="+93" />
                    <RELAYPOSITION athleteid="27512" number="3" reactiontime="+73" />
                    <RELAYPOSITION athleteid="27542" number="4" reactiontime="+91" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="34" agetotalmin="18" gender="X" name="TC Heilbronn 1 GA" number="1">
              <RESULTS>
                <RESULT eventid="1210" reactiontime="+95" swimtime="00:01:12.48" resultid="28539" entrytime="00:01:14.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:17.03" />
                    <SPLIT distance="100" swimtime="00:00:36.42" />
                    <SPLIT distance="150" swimtime="00:00:56.04" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="27505" number="1" reactiontime="+95" />
                    <RELAYPOSITION athleteid="27524" number="2" />
                    <RELAYPOSITION athleteid="27536" number="3" />
                    <RELAYPOSITION athleteid="27507" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
          <OFFICIALS>
            <OFFICIAL officialid="23070" firstname="Udo" gender="M" grade="Tijdwaarnemer" lastname="Schillmüller" nation="GER" />
            <OFFICIAL officialid="27674" firstname="Volker" gender="M" grade="Tijdwaarnemer" lastname="Fabriz" nation="GER" />
            <OFFICIAL officialid="24196" firstname="Marion" gender="F" grade="Team Captain" lastname="Wagner" nation="GER" />
          </OFFICIALS>
        </CLUB>
        <CLUB type="CLUB" code="OCEANUS" nation="NED" clubid="16586" name="Oceanus" shortname="OCEANUS">
          <ATHLETES>
            <ATHLETE firstname="Yvanka" lastname="Ashby" birthdate="2000-04-09" gender="F" nation="NED" license="9020068" athleteid="28450">
              <RESULTS>
                <RESULT eventid="1053" points="407" reactiontime="+123" swimtime="00:00:26.93" resultid="28451" entrytime="00:00:26.83" entrycourse="LCM" />
                <RESULT eventid="1093" points="562" reactiontime="+127" swimtime="00:18:15.33" resultid="28452" entrytime="00:18:55.56" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.47" />
                    <SPLIT distance="100" swimtime="00:01:05.44" />
                    <SPLIT distance="150" swimtime="00:01:40.54" />
                    <SPLIT distance="200" swimtime="00:02:17.19" />
                    <SPLIT distance="250" swimtime="00:02:53.43" />
                    <SPLIT distance="300" swimtime="00:03:29.97" />
                    <SPLIT distance="350" swimtime="00:04:06.32" />
                    <SPLIT distance="400" swimtime="00:04:43.19" />
                    <SPLIT distance="450" swimtime="00:05:19.44" />
                    <SPLIT distance="500" swimtime="00:05:55.98" />
                    <SPLIT distance="550" swimtime="00:06:32.23" />
                    <SPLIT distance="600" swimtime="00:07:08.81" />
                    <SPLIT distance="650" swimtime="00:07:45.29" />
                    <SPLIT distance="700" swimtime="00:08:22.69" />
                    <SPLIT distance="750" swimtime="00:08:59.97" />
                    <SPLIT distance="800" swimtime="00:09:37.30" />
                    <SPLIT distance="850" swimtime="00:10:14.28" />
                    <SPLIT distance="900" swimtime="00:10:51.43" />
                    <SPLIT distance="950" swimtime="00:11:29.22" />
                    <SPLIT distance="1000" swimtime="00:12:06.57" />
                    <SPLIT distance="1050" swimtime="00:12:43.51" />
                    <SPLIT distance="1100" swimtime="00:13:21.44" />
                    <SPLIT distance="1150" swimtime="00:13:59.31" />
                    <SPLIT distance="1200" swimtime="00:14:36.37" />
                    <SPLIT distance="1250" swimtime="00:15:14.05" />
                    <SPLIT distance="1300" swimtime="00:15:51.07" />
                    <SPLIT distance="1350" swimtime="00:16:28.90" />
                    <SPLIT distance="1400" swimtime="00:17:07.74" />
                    <SPLIT distance="1450" swimtime="00:17:43.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1120" points="523" reactiontime="+103" swimtime="00:00:28.94" resultid="28453" entrytime="00:00:30.02" entrycourse="LCM" />
                <RESULT eventid="7278" points="640" reactiontime="+120" swimtime="00:04:19.96" resultid="28454" entrytime="00:04:31.61" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.56" />
                    <SPLIT distance="100" swimtime="00:01:01.13" />
                    <SPLIT distance="150" swimtime="00:01:34.55" />
                    <SPLIT distance="200" swimtime="00:02:08.41" />
                    <SPLIT distance="250" swimtime="00:02:42.15" />
                    <SPLIT distance="300" swimtime="00:03:15.91" />
                    <SPLIT distance="350" swimtime="00:03:49.55" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="C1 - Niet de gehele afstand met het gezicht onder water afgelegd" eventid="1147" reactiontime="+134" status="DSQ" swimtime="00:00:25.09" resultid="28455" />
                <RESULT eventid="1158" points="541" reactiontime="+120" swimtime="00:09:34.58" resultid="28456" entrytime="00:09:18.37" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.25" />
                    <SPLIT distance="100" swimtime="00:01:05.37" />
                    <SPLIT distance="150" swimtime="00:01:40.72" />
                    <SPLIT distance="200" swimtime="00:02:17.38" />
                    <SPLIT distance="250" swimtime="00:02:54.04" />
                    <SPLIT distance="300" swimtime="00:03:31.18" />
                    <SPLIT distance="350" swimtime="00:04:07.95" />
                    <SPLIT distance="400" swimtime="00:04:45.12" />
                    <SPLIT distance="450" swimtime="00:05:22.15" />
                    <SPLIT distance="500" swimtime="00:05:59.21" />
                    <SPLIT distance="550" swimtime="00:06:35.69" />
                    <SPLIT distance="600" swimtime="00:07:13.21" />
                    <SPLIT distance="650" swimtime="00:07:50.24" />
                    <SPLIT distance="700" swimtime="00:08:27.26" />
                    <SPLIT distance="750" swimtime="00:09:02.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="7287" points="520" reactiontime="+123" swimtime="00:00:57.07" resultid="28457" entrytime="00:00:58.52" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1168" points="612" reactiontime="+104" swimtime="00:00:59.84" resultid="28458" entrytime="00:01:01.28" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.69" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ella-May" lastname="Meeuwisse" birthdate="2008-07-21" gender="F" nation="NED" license="9263603" athleteid="28467">
              <RESULTS>
                <RESULT eventid="1147" points="423" reactiontime="+103" swimtime="00:00:25.58" resultid="28468" />
                <RESULT eventid="1168" points="797" reactiontime="+104" swimtime="00:01:01.15" resultid="28469" entrytime="00:01:01.80" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="7287" points="416" reactiontime="+107" swimtime="00:01:03.28" resultid="28470" entrytime="00:01:01.49" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.05" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="100 meter backup" eventid="24851" points="308" reactiontime="+101" swimtime="00:02:36.91" resultid="28471" entrytime="00:02:41.87">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.27" />
                    <SPLIT distance="100" swimtime="00:01:11.58" />
                    <SPLIT distance="150" swimtime="00:01:56.35" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Liam" lastname="Glebbeek" birthdate="1998-01-04" gender="M" nation="NED" license="9010316" athleteid="28459">
              <RESULTS>
                <RESULT eventid="1079" points="528" reactiontime="+96" swimtime="00:00:20.97" resultid="28460" entrytime="00:00:20.54" entrycourse="LCM" />
                <RESULT eventid="7271" points="638" reactiontime="+93" swimtime="00:02:06.57" resultid="28461">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.48" />
                    <SPLIT distance="100" swimtime="00:00:58.76" />
                    <SPLIT distance="150" swimtime="00:01:32.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1127" points="652" reactiontime="+96" swimtime="00:00:23.29" resultid="28462" entrytime="00:00:24.29" entrycourse="LCM" />
                <RESULT eventid="1153" points="639" reactiontime="+115" swimtime="00:00:18.35" resultid="28463" entrytime="00:00:19.28" entrycourse="LCM" />
                <RESULT eventid="1175" points="689" reactiontime="+97" swimtime="00:00:52.25" resultid="28464" entrytime="00:00:51.18">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="7295" points="630" reactiontime="+107" swimtime="00:00:45.96" resultid="28465" entrytime="00:00:52.32" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:21.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1190" points="556" reactiontime="+120" swimtime="00:00:44.43" resultid="28466" entrytime="00:00:45.94">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:21.67" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <OFFICIALS>
            <OFFICIAL officialid="7086" firstname="Ronald" gender="M" grade="Keerpuntcommissaris" lastname="Ashby" nation="NED" />
            <OFFICIAL officialid="25527" firstname="Margret" gender="F" grade="Tijdwaarnemer" lastname="Ashby" nation="NED" />
            <OFFICIAL officialid="6659" firstname="Laura" gender="F" grade="Speaker" lastname="Reemst" nation="NED" />
            <OFFICIAL officialid="6969" firstname="Nico" gender="M" grade="Keerpuntcommissaris" lastname="Langenraad" nameprefix="van" nation="NED" />
            <OFFICIAL officialid="7084" firstname="Owen" gender="M" grade="Tijdwaarnemer" lastname="Ashby" nation="NED" />
            <OFFICIAL officialid="21313" firstname="Nico" gender="M" grade="toezichthouder" lastname="Langeraad" nameprefix="van" nation="NED" />
            <OFFICIAL officialid="6383" firstname="Karin" gender="F" grade="Ploegleider" lastname="Oostveen" nation="NED" />
            <OFFICIAL officialid="2781" firstname="Cassey" gender="F" grade="Tijdwaarnemer" lastname="Glebbeek" nation="NED" />
          </OFFICIALS>
        </CLUB>
        <CLUB type="CLUB" code="TC NEMO" nation="GER" clubid="29262" name="Tauchclub NEMO Plauen e.V." shortname="TC NEMO">
          <ATHLETES>
            <ATHLETE firstname="Hannah" lastname="Troppschuh" birthdate="2009-01-22" gender="F" nation="GER" license="154114000630" athleteid="29263">
              <RESULTS>
                <RESULT eventid="1053" points="1064" reactiontime="+100" swimtime="00:00:20.98" resultid="29264" entrytime="00:00:20.93" />
                <RESULT eventid="1105" points="1445" reactiontime="+121" swimtime="00:03:42.31" resultid="29265" entrytime="00:03:38.74">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:22.87" />
                    <SPLIT distance="100" swimtime="00:00:48.25" />
                    <SPLIT distance="150" swimtime="00:01:15.59" />
                    <SPLIT distance="200" swimtime="00:01:44.54" />
                    <SPLIT distance="250" swimtime="00:02:14.32" />
                    <SPLIT distance="300" swimtime="00:02:43.87" />
                    <SPLIT distance="350" swimtime="00:03:14.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1147" points="961" reactiontime="+105" swimtime="00:00:19.46" resultid="29266" entrytime="00:00:18.78" />
                <RESULT eventid="1182" points="1024" reactiontime="+123" swimtime="00:00:45.12" resultid="29267" entrytime="00:00:43.91">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:21.98" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lotte" lastname="Troppschuh" birthdate="2012-08-18" gender="F" nation="GER" license="15411000631" athleteid="29268">
              <RESULTS>
                <RESULT eventid="1053" points="1498" reactiontime="+97" swimtime="00:00:22.44" resultid="29269" entrytime="00:00:23.28" />
                <RESULT eventid="7278" points="1609" reactiontime="+117" swimtime="00:04:21.81" resultid="29270" entrytime="00:04:34.81">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.38" />
                    <SPLIT distance="100" swimtime="00:01:00.22" />
                    <SPLIT distance="150" swimtime="00:01:33.26" />
                    <SPLIT distance="200" swimtime="00:02:06.75" />
                    <SPLIT distance="250" swimtime="00:02:42.09" />
                    <SPLIT distance="300" swimtime="00:03:16.82" />
                    <SPLIT distance="350" swimtime="00:03:51.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="7287" points="1605" reactiontime="+93" swimtime="00:00:50.37" resultid="29271" entrytime="00:00:51.61">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:23.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="24851" points="1230" reactiontime="+98" swimtime="00:02:03.37" resultid="29272" entrytime="00:02:07.56">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.50" />
                    <SPLIT distance="100" swimtime="00:00:58.69" />
                    <SPLIT distance="150" swimtime="00:01:34.45" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <OFFICIALS>
            <OFFICIAL officialid="27686" firstname="Anne" gender="F" grade="Team Captain" lastname="Lüth" nation="GER" />
          </OFFICIALS>
        </CLUB>
        <CLUB type="CLUB" code="FFESSM" nation="FRA" clubid="22766" name="Team FFESSM France">
          <OFFICIALS>
            <OFFICIAL officialid="24418" firstname="Clément" gender="M" grade="Team Captain" lastname="Normani" nation="FRA" />
          </OFFICIALS>
        </CLUB>
        <CLUB type="CLUB" code="USCO" nation="GER" clubid="22869" name="Unterwasser Sport Club Obertshausen" shortname="Unterwasser Sport Club Obertsh">
          <OFFICIALS>
            <OFFICIAL officialid="24192" firstname="Olha" gender="F" grade="Team Captain" lastname="Zehetbauer" nation="GER" />
          </OFFICIALS>
        </CLUB>
        <CLUB type="CLUB" code="NAUTILUS" nation="BEL" clubid="27608" name="Nautilus Hasselt" shortname="Nautilus" shortname.en="Nautilus Hasselt">
          <ATHLETES>
            <ATHLETE firstname="Mirte" lastname="S&apos;heeren" birthdate="2006-01-01" gender="F" nation="BEL" license="BELF00NAP011381" athleteid="29146">
              <RESULTS>
                <RESULT eventid="7254" points="832" reactiontime="+90" swimtime="00:02:06.93" resultid="29164" entrytime="00:01:57.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.57" />
                    <SPLIT distance="100" swimtime="00:01:02.20" />
                    <SPLIT distance="150" swimtime="00:01:35.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1120" points="815" reactiontime="+88" swimtime="00:00:25.84" resultid="29165" entrytime="00:00:25.00" />
                <RESULT eventid="1168" points="757" reactiontime="+90" swimtime="00:00:58.35" resultid="29166" entrytime="00:00:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.34" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Stijn" lastname="Maes" birthdate="1992-01-01" gender="M" nation="BEL" license="BELF00NAP000144" athleteid="27641">
              <RESULTS>
                <RESULT eventid="16574" points="378" reactiontime="+96" swimtime="00:09:30.93" resultid="29170" entrytime="00:10:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.98" />
                    <SPLIT distance="100" swimtime="00:00:58.44" />
                    <SPLIT distance="150" swimtime="00:01:32.82" />
                    <SPLIT distance="200" swimtime="00:02:09.15" />
                    <SPLIT distance="250" swimtime="00:02:45.69" />
                    <SPLIT distance="300" swimtime="00:03:22.32" />
                    <SPLIT distance="350" swimtime="00:03:59.26" />
                    <SPLIT distance="400" swimtime="00:04:36.31" />
                    <SPLIT distance="450" swimtime="00:05:13.21" />
                    <SPLIT distance="500" swimtime="00:05:50.88" />
                    <SPLIT distance="550" swimtime="00:06:28.53" />
                    <SPLIT distance="600" swimtime="00:07:06.33" />
                    <SPLIT distance="650" swimtime="00:07:43.73" />
                    <SPLIT distance="700" swimtime="00:08:22.22" />
                    <SPLIT distance="750" swimtime="00:08:56.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1203" points="604" reactiontime="+103" swimtime="00:04:30.67" resultid="29171" entrytime="00:04:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.37" />
                    <SPLIT distance="100" swimtime="00:00:59.84" />
                    <SPLIT distance="150" swimtime="00:01:33.47" />
                    <SPLIT distance="200" swimtime="00:02:08.39" />
                    <SPLIT distance="250" swimtime="00:02:44.40" />
                    <SPLIT distance="300" swimtime="00:03:20.84" />
                    <SPLIT distance="350" swimtime="00:03:56.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="18215" points="425" reactiontime="+104" swimtime="00:17:48.64" resultid="29462" entrytime="00:18:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.90" />
                    <SPLIT distance="100" swimtime="00:00:58.82" />
                    <SPLIT distance="150" swimtime="00:01:32.10" />
                    <SPLIT distance="200" swimtime="00:02:07.35" />
                    <SPLIT distance="250" swimtime="00:02:43.51" />
                    <SPLIT distance="300" swimtime="00:03:19.92" />
                    <SPLIT distance="350" swimtime="00:03:56.02" />
                    <SPLIT distance="400" swimtime="00:04:32.15" />
                    <SPLIT distance="450" swimtime="00:05:08.78" />
                    <SPLIT distance="500" swimtime="00:05:45.97" />
                    <SPLIT distance="550" swimtime="00:06:22.03" />
                    <SPLIT distance="600" swimtime="00:06:59.37" />
                    <SPLIT distance="650" swimtime="00:07:35.72" />
                    <SPLIT distance="700" swimtime="00:08:13.29" />
                    <SPLIT distance="750" swimtime="00:08:50.03" />
                    <SPLIT distance="800" swimtime="00:09:25.57" />
                    <SPLIT distance="850" swimtime="00:10:01.44" />
                    <SPLIT distance="900" swimtime="00:10:37.74" />
                    <SPLIT distance="950" swimtime="00:11:13.99" />
                    <SPLIT distance="1000" swimtime="00:11:51.23" />
                    <SPLIT distance="1050" swimtime="00:12:27.28" />
                    <SPLIT distance="1100" swimtime="00:13:03.94" />
                    <SPLIT distance="1150" swimtime="00:13:40.80" />
                    <SPLIT distance="1200" swimtime="00:14:17.20" />
                    <SPLIT distance="1250" swimtime="00:14:53.48" />
                    <SPLIT distance="1300" swimtime="00:15:29.73" />
                    <SPLIT distance="1350" swimtime="00:16:05.49" />
                    <SPLIT distance="1400" swimtime="00:16:41.90" />
                    <SPLIT distance="1450" swimtime="00:17:14.41" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Koen" lastname="Merken" birthdate="1989-01-01" gender="M" nation="BEL" license="NELOS 47020" athleteid="29149">
              <RESULTS>
                <RESULT eventid="7271" points="637" reactiontime="+97" swimtime="00:02:06.61" resultid="29162" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.45" />
                    <SPLIT distance="100" swimtime="00:00:59.65" />
                    <SPLIT distance="150" swimtime="00:01:32.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1127" points="461" reactiontime="+91" swimtime="00:00:26.13" resultid="29163" entrytime="00:00:26.85" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Wouter" lastname="Rabijns" birthdate="1990-01-01" gender="M" nation="BEL" license="BELF00NAP011380" athleteid="29148">
              <RESULTS>
                <RESULT eventid="7271" points="762" reactiontime="+99" swimtime="00:01:59.27" resultid="29172" entrytime="00:01:54.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.34" />
                    <SPLIT distance="100" swimtime="00:00:56.11" />
                    <SPLIT distance="150" swimtime="00:01:27.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1127" points="548" reactiontime="+102" swimtime="00:00:24.67" resultid="29173" entrytime="00:00:24.96" />
                <RESULT eventid="1175" points="618" reactiontime="+102" swimtime="00:00:54.19" resultid="29174" entrytime="00:00:54.70">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1203" points="711" reactiontime="+104" swimtime="00:04:16.38" resultid="29175" entrytime="00:04:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.39" />
                    <SPLIT distance="100" swimtime="00:00:59.73" />
                    <SPLIT distance="150" swimtime="00:01:32.40" />
                    <SPLIT distance="200" swimtime="00:02:05.95" />
                    <SPLIT distance="250" swimtime="00:02:39.30" />
                    <SPLIT distance="300" swimtime="00:03:12.64" />
                    <SPLIT distance="350" swimtime="00:03:45.52" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Elise" lastname="Croes" birthdate="2004-01-01" gender="F" nation="BEL" license="BELF00NAP011365" athleteid="27634">
              <RESULTS>
                <RESULT eventid="7254" points="1015" reactiontime="+82" swimtime="00:01:49.98" resultid="29150" entrytime="00:01:51.79">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.76" />
                    <SPLIT distance="100" swimtime="00:00:53.90" />
                    <SPLIT distance="150" swimtime="00:01:22.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1120" points="997" reactiontime="+85" swimtime="00:00:23.35" resultid="29151" entrytime="00:00:23.10" />
                <RESULT eventid="1168" points="1020" reactiontime="+85" swimtime="00:00:50.46" resultid="29152" entrytime="00:00:51.18">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:24.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1196" points="1396" reactiontime="+86" swimtime="00:03:56.28" resultid="29153" entrytime="00:03:57.28">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.03" />
                    <SPLIT distance="100" swimtime="00:00:56.69" />
                    <SPLIT distance="150" swimtime="00:01:26.98" />
                    <SPLIT distance="200" swimtime="00:01:57.33" />
                    <SPLIT distance="250" swimtime="00:02:27.17" />
                    <SPLIT distance="300" swimtime="00:02:57.38" />
                    <SPLIT distance="350" swimtime="00:03:27.48" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Linda" lastname="Quintiens" birthdate="1963-01-01" gender="F" nation="BEL" license="BELF00NAP011377" athleteid="27644">
              <RESULTS>
                <RESULT eventid="7254" points="8058" reactiontime="+109" swimtime="00:02:59.56" resultid="29158" entrytime="00:02:51.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.18" />
                    <SPLIT distance="100" swimtime="00:01:25.16" />
                    <SPLIT distance="150" swimtime="00:02:13.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1120" points="626" reactiontime="+105" swimtime="00:00:36.26" resultid="29159" entrytime="00:00:36.92" />
                <RESULT eventid="1168" points="580" reactiontime="+104" swimtime="00:01:19.68" resultid="29160" entrytime="00:01:21.60">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1196" points="4413" reactiontime="+109" swimtime="00:06:05.78" resultid="29161" entrytime="00:06:07.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.04" />
                    <SPLIT distance="100" swimtime="00:01:24.52" />
                    <SPLIT distance="150" swimtime="00:02:11.90" />
                    <SPLIT distance="200" swimtime="00:02:59.77" />
                    <SPLIT distance="250" swimtime="00:03:47.45" />
                    <SPLIT distance="300" swimtime="00:04:35.09" />
                    <SPLIT distance="350" swimtime="00:05:21.35" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="René" lastname="Hendrikx" birthdate="1993-01-01" gender="M" nation="BEL" license="BELF00NAP011376" athleteid="27638">
              <RESULTS>
                <RESULT eventid="1175" points="503" reactiontime="+97" swimtime="00:00:58.01" resultid="29167" entrytime="00:00:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1203" points="513" reactiontime="+99" swimtime="00:04:45.80" resultid="29168" entrytime="00:04:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.08" />
                    <SPLIT distance="100" swimtime="00:01:03.33" />
                    <SPLIT distance="150" swimtime="00:01:38.49" />
                    <SPLIT distance="200" swimtime="00:02:15.00" />
                    <SPLIT distance="250" swimtime="00:02:52.53" />
                    <SPLIT distance="300" swimtime="00:03:30.78" />
                    <SPLIT distance="350" swimtime="00:04:08.70" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Hasan" lastname="Eryilmaz" birthdate="2008-01-01" gender="M" nation="BEL" license="NELOS 50217" athleteid="29147">
              <RESULTS>
                <RESULT eventid="7271" points="858" reactiontime="+91" swimtime="00:01:59.34" resultid="29154" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.96" />
                    <SPLIT distance="100" swimtime="00:00:55.85" />
                    <SPLIT distance="150" swimtime="00:01:27.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1127" points="820" reactiontime="+87" swimtime="00:00:24.43" resultid="29155" entrytime="00:00:25.00" />
                <RESULT eventid="1153" status="WDR" swimtime="00:00:00.00" resultid="29156" entrytime="00:00:24.00" />
                <RESULT eventid="1175" status="WDR" swimtime="00:00:00.00" resultid="29157" entrytime="00:00:57.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="34" agemin="18" agetotalmax="-1" agetotalmin="-1" gender="X" name="Team Nautilus GA" number="1">
              <RESULTS>
                <RESULT eventid="1140" reactiontime="+84" swimtime="00:03:37.56" resultid="29176" entrytime="00:04:31.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:24.85" />
                    <SPLIT distance="100" swimtime="00:00:50.89" />
                    <SPLIT distance="150" swimtime="00:01:17.94" />
                    <SPLIT distance="200" swimtime="00:01:47.87" />
                    <SPLIT distance="250" swimtime="00:02:14.26" />
                    <SPLIT distance="300" swimtime="00:02:42.53" />
                    <SPLIT distance="350" swimtime="00:03:08.32" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="27634" number="1" reactiontime="+84" />
                    <RELAYPOSITION athleteid="29146" number="2" reactiontime="+57" />
                    <RELAYPOSITION athleteid="29148" number="3" reactiontime="+72" />
                    <RELAYPOSITION athleteid="27641" number="4" reactiontime="+61" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="34" agetotalmin="18" gender="X" name="Team Nautilus GA" number="1">
              <RESULTS>
                <RESULT comment="Backup 50 meter" eventid="1210" reactiontime="+89" swimtime="00:01:45.55" resultid="29177" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:19.18" />
                    <SPLIT distance="100" swimtime="00:00:46.08" />
                    <SPLIT distance="150" swimtime="00:01:14.86" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="27634" number="1" reactiontime="+89" />
                    <RELAYPOSITION athleteid="29146" number="2" reactiontime="+35" />
                    <RELAYPOSITION athleteid="29148" number="3" reactiontime="+100" />
                    <RELAYPOSITION athleteid="27641" number="4" reactiontime="+62" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
          <COACHES>
            <COACH firstname="Free" gender="M" lastname="Deurinckx" nation="BEL" type="COACH" />
          </COACHES>
          <OFFICIALS>
            <OFFICIAL officialid="24573" firstname="Stijn" gender="M" grade="Team Captain" lastname="Maes" nation="BEL" />
            <OFFICIAL officialid="24080" firstname="Free" gender="M" grade="Lijnrechter" lastname="Duerinckx" nation="BEL" />
          </OFFICIALS>
        </CLUB>
        <CLUB type="CLUB" code="SGD" nation="GER" clubid="22402" name="SG Dresden">
          <COACHES>
            <COACH firstname="Sven" gender="M" lastname="Klabunde" nation="GER" />
          </COACHES>
          <OFFICIALS>
            <OFFICIAL officialid="26165" firstname="Sven" gender="M" grade="Team Captain" lastname="Klabunde" nation="GER" />
          </OFFICIALS>
        </CLUB>
        <CLUB type="CLUB" code="VZ UTRECHT" nation="NED" clubid="18179" name="Vinzwemmen Utrecht" shortname="VZ Utrecht">
          <ATHLETES>
            <ATHLETE firstname="Niels" lastname="van den Brom" birthdate="1989-03-05" gender="M" nation="NED" license="9265749" athleteid="29368">
              <RESULTS>
                <RESULT eventid="1079" points="334" reactiontime="+92" swimtime="00:00:24.42" resultid="29369" entrytime="00:00:24.52" entrycourse="LCM" />
                <RESULT eventid="7271" points="501" reactiontime="+90" swimtime="00:02:17.13" resultid="29370">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.53" />
                    <SPLIT distance="100" swimtime="00:01:05.51" />
                    <SPLIT distance="150" swimtime="00:01:41.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1127" points="487" reactiontime="+98" swimtime="00:00:25.66" resultid="29371" />
                <RESULT eventid="1153" points="304" reactiontime="+106" swimtime="00:00:23.51" resultid="29372" />
                <RESULT eventid="1175" points="517" reactiontime="+94" swimtime="00:00:57.49" resultid="29373" entrytime="00:00:58.77" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="24862" points="352" reactiontime="+112" swimtime="00:02:10.17" resultid="29374">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.59" />
                    <SPLIT distance="100" swimtime="00:01:02.27" />
                    <SPLIT distance="150" swimtime="00:01:36.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="7295" points="332" reactiontime="+99" swimtime="00:00:56.89" resultid="29375" entrytime="00:00:57.66" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.30" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Brian" lastname="Joosten" birthdate="1972-12-24" gender="M" nation="NED" license="34212" athleteid="29350">
              <RESULTS>
                <RESULT comment="Nederlands Record, Nederlands record" eventid="1079" points="1080" reactiontime="+98" swimtime="00:00:20.72" resultid="29351" entrytime="00:00:21.26" entrycourse="LCM" />
                <RESULT comment="Nederlands record" eventid="7271" points="1017" reactiontime="+99" swimtime="00:01:56.93" resultid="29352" entrytime="00:01:57.59" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.05" />
                    <SPLIT distance="100" swimtime="00:00:56.58" />
                    <SPLIT distance="150" swimtime="00:01:26.97" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Nederlands record" eventid="1127" points="902" reactiontime="+101" swimtime="00:00:23.69" resultid="29353" entrytime="00:00:23.89" entrycourse="LCM" />
                <RESULT comment="Nederlands record" eventid="1153" points="1045" reactiontime="+98" swimtime="00:00:18.25" resultid="29354" entrytime="00:00:18.38" entrycourse="LCM" />
                <RESULT comment="Nederlands record" eventid="1175" points="1017" reactiontime="+98" swimtime="00:00:51.60" resultid="29355" entrytime="00:00:51.90" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:24.91" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Nederlands record" eventid="7295" points="1050" reactiontime="+102" swimtime="00:00:47.47" resultid="29356" entrytime="00:00:48.25" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:23.03" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Nederlands record" eventid="1190" points="1142" reactiontime="+138" swimtime="00:00:45.37" resultid="29357" entrytime="00:00:48.10" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:21.66" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Nederlands record" eventid="24862" points="1038" reactiontime="+115" swimtime="00:01:51.37" resultid="29358" entrytime="00:01:45.81" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.18" />
                    <SPLIT distance="100" swimtime="00:00:55.33" />
                    <SPLIT distance="150" swimtime="00:01:25.62" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Zoë" lastname="Bommel" birthdate="2013-07-13" gender="F" nation="NED" license="9263554" athleteid="29279">
              <RESULTS>
                <RESULT eventid="1053" points="520" reactiontime="+95" swimtime="00:00:31.92" resultid="29280" entrytime="00:00:31.54" entrycourse="LCM" />
                <RESULT eventid="1120" points="570" reactiontime="+104" swimtime="00:00:36.03" resultid="29281" entrytime="00:00:35.54" entrycourse="LCM" />
                <RESULT eventid="1168" points="567" reactiontime="+99" swimtime="00:01:17.94" resultid="29282" entrytime="00:01:19.27" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="7287" points="502" reactiontime="+106" swimtime="00:01:14.17" resultid="29283" entrytime="00:01:15.93" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="24851" points="484" reactiontime="+118" swimtime="00:02:48.34" resultid="29284" entrytime="00:02:49.66" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.12" />
                    <SPLIT distance="100" swimtime="00:01:21.26" />
                    <SPLIT distance="150" swimtime="00:02:06.64" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lars" lastname="Jong" birthdate="2010-04-10" gender="M" nameprefix="de" nation="NED" license="9265751" athleteid="29335">
              <RESULTS>
                <RESULT eventid="1079" points="733" reactiontime="+94" swimtime="00:00:26.13" resultid="29336" entrytime="00:00:28.57" />
                <RESULT eventid="7271" points="843" reactiontime="+103" swimtime="00:02:27.67" resultid="29337">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.57" />
                    <SPLIT distance="100" swimtime="00:01:09.19" />
                    <SPLIT distance="150" swimtime="00:01:49.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1127" points="908" reactiontime="+97" swimtime="00:00:27.58" resultid="29338" entrytime="00:00:30.21" />
                <RESULT eventid="1175" points="687" reactiontime="+88" swimtime="00:01:03.86" resultid="29339" entrytime="00:01:07.40">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="7295" points="748" reactiontime="+88" swimtime="00:00:59.97" resultid="29340" entrytime="00:01:09.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="24862" points="656" reactiontime="+96" swimtime="00:02:19.06" resultid="29341" entrytime="00:02:45.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.50" />
                    <SPLIT distance="100" swimtime="00:01:07.61" />
                    <SPLIT distance="150" swimtime="00:01:47.06" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Erik" lastname="Jong" birthdate="1969-02-03" gender="M" nameprefix="de" nation="NED" license="9036495" athleteid="29328">
              <RESULTS>
                <RESULT eventid="1079" points="684" reactiontime="+107" swimtime="00:00:24.12" resultid="29329" entrytime="00:00:24.65" entrycourse="LCM" />
                <RESULT eventid="7271" points="761" reactiontime="+103" swimtime="00:02:08.77" resultid="29330" entrytime="00:02:09.04" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.70" />
                    <SPLIT distance="100" swimtime="00:01:01.75" />
                    <SPLIT distance="150" swimtime="00:01:35.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="7264" points="699" reactiontime="+112" swimtime="00:04:31.39" resultid="29331" entrytime="00:04:29.46" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.51" />
                    <SPLIT distance="100" swimtime="00:01:05.61" />
                    <SPLIT distance="150" swimtime="00:01:39.37" />
                    <SPLIT distance="200" swimtime="00:02:13.61" />
                    <SPLIT distance="250" swimtime="00:02:48.22" />
                    <SPLIT distance="300" swimtime="00:03:23.89" />
                    <SPLIT distance="350" swimtime="00:03:58.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1153" points="696" reactiontime="+99" swimtime="00:00:20.89" resultid="29332" entrytime="00:00:20.83" entrycourse="LCM" />
                <RESULT eventid="1203" points="970" reactiontime="+108" swimtime="00:04:47.75" resultid="29333" entrytime="00:04:42.63" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.24" />
                    <SPLIT distance="100" swimtime="00:01:03.74" />
                    <SPLIT distance="150" swimtime="00:01:38.63" />
                    <SPLIT distance="200" swimtime="00:02:15.54" />
                    <SPLIT distance="250" swimtime="00:02:53.24" />
                    <SPLIT distance="300" swimtime="00:03:31.31" />
                    <SPLIT distance="350" swimtime="00:04:10.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="24862" points="708" reactiontime="+114" swimtime="00:02:06.49" resultid="29334" entrytime="00:02:04.38" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.25" />
                    <SPLIT distance="100" swimtime="00:01:00.97" />
                    <SPLIT distance="150" swimtime="00:01:34.26" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Aizza" lastname="Bommel" birthdate="2011-12-14" gender="F" nation="NED" license="9263553" athleteid="29273">
              <RESULTS>
                <RESULT comment="A1 - Bewogen of te vroeg weg bij de start (geen tijd noteren)" eventid="1053" reactiontime="+52" status="DSQ" swimtime="00:00:00.00" resultid="29274" entrytime="00:00:31.77" entrycourse="LCM" />
                <RESULT eventid="1120" points="547" swimtime="00:00:33.37" resultid="29275" entrytime="00:00:33.14" entrycourse="LCM" />
                <RESULT eventid="1168" points="441" reactiontime="+77" swimtime="00:01:17.69" resultid="29276" entrytime="00:01:20.06" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="7287" points="343" reactiontime="+67" swimtime="00:01:11.73" resultid="29277" entrytime="00:01:13.78" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.51" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="A1 - Bewogen of te vroeg weg bij de start (geen tijd noteren)" eventid="24851" reactiontime="+51" status="DSQ" swimtime="00:02:43.28" resultid="29278" entrytime="00:02:49.44" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.04" />
                    <SPLIT distance="100" swimtime="00:01:18.75" />
                    <SPLIT distance="150" swimtime="00:02:03.57" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Nikolai" lastname="Kanin" birthdate="2013-10-23" gender="M" nation="RUS" license="9265752" athleteid="29359">
              <RESULTS>
                <RESULT eventid="1079" points="595" reactiontime="+109" swimtime="00:00:33.00" resultid="29360" entrytime="00:00:34.35" entrycourse="LCM" />
                <RESULT eventid="1127" points="541" swimtime="00:00:36.91" resultid="29361" entrytime="00:00:39.23" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Laura" lastname="Spanjers" birthdate="1993-08-04" gender="F" nation="NED" license="9259545" athleteid="29362">
              <RESULTS>
                <RESULT eventid="1053" points="593" reactiontime="+99" swimtime="00:00:23.75" resultid="29363" entrytime="00:00:23.78" entrycourse="LCM" />
                <RESULT eventid="1120" points="675" reactiontime="+92" swimtime="00:00:26.59" resultid="29364" entrytime="00:00:27.27" entrycourse="LCM" />
                <RESULT eventid="1147" points="485" reactiontime="+108" swimtime="00:00:23.98" resultid="29365" entrytime="00:00:22.60" entrycourse="LCM" />
                <RESULT eventid="1168" points="649" reactiontime="+89" swimtime="00:00:58.68" resultid="29366" entrytime="00:00:59.79" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="7287" points="631" reactiontime="+102" swimtime="00:00:53.53" resultid="29367" entrytime="00:00:53.18" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.33" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Hélène" lastname="Bouwmeester" birthdate="1995-04-02" gender="F" nation="NED" license="9218747" athleteid="29297">
              <RESULTS>
                <RESULT eventid="1053" points="583" reactiontime="+105" swimtime="00:00:23.88" resultid="29298" entrytime="00:00:23.01" entrycourse="LCM" />
                <RESULT eventid="7278" points="629" reactiontime="+106" swimtime="00:04:21.53" resultid="29299" entrytime="00:04:14.69" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.40" />
                    <SPLIT distance="100" swimtime="00:01:00.83" />
                    <SPLIT distance="150" swimtime="00:01:34.81" />
                    <SPLIT distance="200" swimtime="00:02:09.31" />
                    <SPLIT distance="250" swimtime="00:02:43.59" />
                    <SPLIT distance="300" swimtime="00:03:17.84" />
                    <SPLIT distance="350" swimtime="00:03:50.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1147" points="624" reactiontime="+94" swimtime="00:00:22.05" resultid="29300" entrytime="00:00:21.60" entrycourse="LCM" />
                <RESULT eventid="7287" points="699" reactiontime="+101" swimtime="00:00:51.74" resultid="29301" entrytime="00:00:51.97" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:24.56" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Hanna" lastname="Bouhuis" birthdate="2001-08-20" gender="F" nation="NED" license="9024271" athleteid="29291">
              <RESULTS>
                <RESULT eventid="1053" points="597" reactiontime="+115" swimtime="00:00:23.70" resultid="29292" entrytime="00:00:24.49" entrycourse="LCM" />
                <RESULT eventid="7278" points="583" reactiontime="+112" swimtime="00:04:28.16" resultid="29293" entrytime="00:04:33.81" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.56" />
                    <SPLIT distance="100" swimtime="00:01:04.19" />
                    <SPLIT distance="150" swimtime="00:01:39.66" />
                    <SPLIT distance="200" swimtime="00:02:15.91" />
                    <SPLIT distance="250" swimtime="00:02:50.30" />
                    <SPLIT distance="300" swimtime="00:03:24.83" />
                    <SPLIT distance="350" swimtime="00:03:58.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1147" status="WDR" swimtime="00:00:00.00" resultid="29294" entrytime="00:00:21.63" entrycourse="LCM" />
                <RESULT eventid="7287" status="WDR" swimtime="00:00:00.00" resultid="29295" entrytime="00:00:58.86" entrycourse="LCM" />
                <RESULT eventid="24851" status="WDR" swimtime="00:00:00.00" resultid="29296" entrytime="00:01:59.51" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lucie" lastname="Gout" birthdate="2012-04-01" gender="F" nation="NED" license="9263557" athleteid="29316">
              <RESULTS>
                <RESULT comment="A1 - Bewogen of te vroeg weg bij de start (geen tijd noteren)" eventid="1053" reactiontime="+69" status="DSQ" swimtime="00:00:34.72" resultid="29317" entrytime="00:00:34.30" entrycourse="LCM" />
                <RESULT eventid="7254" points="749" reactiontime="+117" swimtime="00:02:53.02" resultid="29318">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.46" />
                    <SPLIT distance="100" swimtime="00:01:23.81" />
                    <SPLIT distance="150" swimtime="00:02:11.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1120" points="741" reactiontime="+115" swimtime="00:00:33.02" resultid="29319" entrytime="00:00:35.12" entrycourse="LCM" />
                <RESULT eventid="1168" points="634" reactiontime="+108" swimtime="00:01:15.07" resultid="29320" entrytime="00:01:17.88" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.76" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="geen 50 meter tijd" eventid="7287" points="338" reactiontime="+114" swimtime="00:01:24.60" resultid="29321" entrytime="00:01:22.60" entrycourse="LCM" />
                <RESULT eventid="24851" points="334" reactiontime="+122" swimtime="00:03:10.44" resultid="29322" entrytime="00:03:02.70" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.22" />
                    <SPLIT distance="100" swimtime="00:01:30.83" />
                    <SPLIT distance="150" swimtime="00:02:23.09" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Floor" lastname="Boon" birthdate="2010-06-08" gender="F" nation="NED" license="9255534" athleteid="29285">
              <RESULTS>
                <RESULT eventid="1053" points="1000" reactiontime="+92" swimtime="00:00:22.70" resultid="29286" entrytime="00:00:22.89" entrycourse="LCM" />
                <RESULT comment="Nederlands record" eventid="7278" points="1023" reactiontime="+80" swimtime="00:04:33.80" resultid="29287" entrytime="00:04:45.51" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.68" />
                    <SPLIT distance="100" swimtime="00:01:03.47" />
                    <SPLIT distance="150" swimtime="00:01:38.13" />
                    <SPLIT distance="200" swimtime="00:02:14.32" />
                    <SPLIT distance="250" swimtime="00:02:50.14" />
                    <SPLIT distance="300" swimtime="00:03:25.90" />
                    <SPLIT distance="350" swimtime="00:04:01.36" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Nederlands record" eventid="1168" points="1024" reactiontime="+77" swimtime="00:00:58.68" resultid="29288" entrytime="00:00:58.79" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="7287" points="974" reactiontime="+90" swimtime="00:00:50.66" resultid="29289" entrytime="00:00:51.71" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:23.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="24851" points="1127" reactiontime="+90" swimtime="00:02:00.43" resultid="29290" entrytime="00:01:58.28" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.60" />
                    <SPLIT distance="100" swimtime="00:00:58.53" />
                    <SPLIT distance="150" swimtime="00:01:30.69" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bodijne" lastname="Chaitram" birthdate="2009-09-12" gender="F" nation="NED" license="9263555" athleteid="29302">
              <RESULTS>
                <RESULT eventid="1053" points="369" reactiontime="+89" swimtime="00:00:29.86" resultid="29303" entrytime="00:00:29.02" entrycourse="LCM" />
                <RESULT eventid="7254" points="590" reactiontime="+103" swimtime="00:02:31.07" resultid="29304">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.91" />
                    <SPLIT distance="100" swimtime="00:01:13.74" />
                    <SPLIT distance="150" swimtime="00:01:53.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1120" points="537" reactiontime="+93" swimtime="00:00:30.54" resultid="29305" entrytime="00:00:31.36" entrycourse="LCM" />
                <RESULT eventid="1168" points="564" reactiontime="+103" swimtime="00:01:08.60" resultid="29306" entrytime="00:01:11.18" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="7287" points="298" reactiontime="+92" swimtime="00:01:10.70" resultid="29307" entrytime="00:01:07.26" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="24851" points="286" reactiontime="+98" swimtime="00:02:40.89" resultid="29308" entrytime="00:03:06.33" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.80" />
                    <SPLIT distance="100" swimtime="00:01:15.26" />
                    <SPLIT distance="150" swimtime="00:02:01.53" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Saphine" lastname="Chaitram" birthdate="2011-12-07" gender="F" nation="NED" license="9263556" athleteid="29309">
              <RESULTS>
                <RESULT eventid="1053" points="359" reactiontime="+103" swimtime="00:00:31.92" resultid="29310" entrytime="00:00:32.87" entrycourse="LCM" />
                <RESULT eventid="7254" points="445" reactiontime="+100" swimtime="00:02:56.97" resultid="29311">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.14" />
                    <SPLIT distance="100" swimtime="00:01:29.94" />
                    <SPLIT distance="150" swimtime="00:02:16.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1120" points="442" reactiontime="+103" swimtime="00:00:35.83" resultid="29312" entrytime="00:00:35.18" entrycourse="LCM" />
                <RESULT eventid="1168" points="403" reactiontime="+104" swimtime="00:01:20.02" resultid="29313" entrytime="00:01:22.45" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="7287" points="264" reactiontime="+106" swimtime="00:01:18.26" resultid="29314" entrytime="00:01:19.99" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="24851" points="376" reactiontime="+105" swimtime="00:02:53.55" resultid="29315" entrytime="00:03:04.30" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.90" />
                    <SPLIT distance="100" swimtime="00:01:25.34" />
                    <SPLIT distance="150" swimtime="00:02:12.68" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marije" lastname="Jansen" birthdate="1985-09-29" gender="F" nation="NED" license="9265498" athleteid="29323">
              <RESULTS>
                <RESULT comment="Nederlands record" eventid="1147" points="1248" reactiontime="+94" swimtime="00:00:19.90" resultid="29324" entrytime="00:00:20.41" entrycourse="LCM" />
                <RESULT comment="Nederlands record" eventid="1168" points="1362" reactiontime="+89" swimtime="00:00:54.64" resultid="29325" entrytime="00:00:56.79" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.24" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Nederlands record" eventid="7287" points="1223" reactiontime="+94" swimtime="00:00:50.39" resultid="29326" entrytime="00:00:49.35" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:24.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="24851" points="1120" reactiontime="+95" swimtime="00:01:58.34" resultid="29327" entrytime="00:01:57.39" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.19" />
                    <SPLIT distance="100" swimtime="00:00:56.76" />
                    <SPLIT distance="150" swimtime="00:01:27.73" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Anyk" lastname="Joosten" birthdate="2005-12-01" gender="F" nation="NED" license="9220510" athleteid="29342">
              <RESULTS>
                <RESULT eventid="1053" points="517" reactiontime="+113" swimtime="00:00:24.86" resultid="29343" entrytime="00:00:24.55" entrycourse="LCM" />
                <RESULT eventid="7254" points="536" reactiontime="+92" swimtime="00:02:16.07" resultid="29344" entrytime="00:02:20.04" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.11" />
                    <SPLIT distance="100" swimtime="00:01:03.37" />
                    <SPLIT distance="150" swimtime="00:01:40.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="7278" points="455" reactiontime="+97" swimtime="00:04:51.29" resultid="29345" entrytime="00:04:45.70" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.29" />
                    <SPLIT distance="100" swimtime="00:01:09.18" />
                    <SPLIT distance="150" swimtime="00:01:45.95" />
                    <SPLIT distance="200" swimtime="00:02:23.05" />
                    <SPLIT distance="250" swimtime="00:03:00.61" />
                    <SPLIT distance="300" swimtime="00:03:38.61" />
                    <SPLIT distance="350" swimtime="00:04:16.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1147" points="515" reactiontime="+107" swimtime="00:00:23.51" resultid="29346" entrytime="00:00:22.96" entrycourse="LCM" />
                <RESULT eventid="1168" points="571" reactiontime="+97" swimtime="00:01:01.21" resultid="29347" entrytime="00:01:02.06" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="7287" points="577" reactiontime="+110" swimtime="00:00:55.13" resultid="29348" entrytime="00:00:57.65" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1182" points="390" reactiontime="+118" swimtime="00:01:00.44" resultid="29349">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.76" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="34" agetotalmin="18" gender="M" name="VZU HA" number="3">
              <RESULTS>
                <RESULT comment="E1 - Te vroeg overgenomen, waarna niet teruggekeerd naar de bassinwand om opnieuw te vertrekken, 2e zwemmer te vroeg" eventid="24873" reactiontime="+99" status="DSQ" swimtime="00:00:00.00" resultid="29376" entrytime="00:03:50.71">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.19" />
                    <SPLIT distance="100" swimtime="00:00:57.54" />
                    <SPLIT distance="150" swimtime="00:01:22.83" />
                    <SPLIT distance="200" swimtime="00:01:52.40" />
                    <SPLIT distance="250" swimtime="00:02:20.74" />
                    <SPLIT distance="300" swimtime="00:02:52.14" />
                    <SPLIT distance="350" swimtime="00:03:15.16" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="29368" number="1" reactiontime="+99" status="DSQ" />
                    <RELAYPOSITION athleteid="29328" number="2" reactiontime="-16" status="DSQ" />
                    <RELAYPOSITION athleteid="29335" number="3" reactiontime="+65" status="DSQ" />
                    <RELAYPOSITION athleteid="29350" number="4" reactiontime="+17" status="DSQ" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="34" agetotalmin="18" gender="M" name="VZU HA BM" number="3">
              <RESULTS>
                <RESULT eventid="26768" reactiontime="+100" status="EXH" swimtime="00:01:50.73" resultid="29377" entrytime="00:01:39.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.91" />
                    <SPLIT distance="100" swimtime="00:01:00.05" />
                    <SPLIT distance="150" swimtime="00:01:26.91" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="29368" number="1" reactiontime="+100" />
                    <RELAYPOSITION athleteid="29359" number="2" reactiontime="+31" />
                    <RELAYPOSITION athleteid="29335" number="3" reactiontime="+53" />
                    <RELAYPOSITION athleteid="29328" number="4" reactiontime="+24" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="34" agetotalmin="18" gender="F" name="VZU DA" number="1">
              <RESULTS>
                <RESULT eventid="1217" reactiontime="+98" swimtime="00:03:28.41" resultid="29378" entrytime="00:03:32.63">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:24.83" />
                    <SPLIT distance="100" swimtime="00:00:51.49" />
                    <SPLIT distance="150" swimtime="00:01:16.09" />
                    <SPLIT distance="200" swimtime="00:01:43.75" />
                    <SPLIT distance="250" swimtime="00:02:09.43" />
                    <SPLIT distance="300" swimtime="00:02:37.59" />
                    <SPLIT distance="350" swimtime="00:03:01.60" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="29323" number="1" reactiontime="+98" />
                    <RELAYPOSITION athleteid="29297" number="2" reactiontime="+37" />
                    <RELAYPOSITION athleteid="29362" number="3" reactiontime="+33" />
                    <RELAYPOSITION athleteid="29285" number="4" reactiontime="+47" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="34" agetotalmin="18" gender="F" name="VZU DA" number="1">
              <RESULTS>
                <RESULT comment="Nederlands record" eventid="26758" reactiontime="+99" swimtime="00:01:34.01" resultid="29379" entrytime="00:01:33.34">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:23.65" />
                    <SPLIT distance="100" swimtime="00:00:48.02" />
                    <SPLIT distance="150" swimtime="00:01:11.55" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="29297" number="1" reactiontime="+99" />
                    <RELAYPOSITION athleteid="29342" number="2" reactiontime="+26" />
                    <RELAYPOSITION athleteid="29362" number="3" reactiontime="+17" />
                    <RELAYPOSITION athleteid="29285" number="4" reactiontime="+32" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="13" agemin="12" agetotalmax="-1" agetotalmin="-1" gender="F" name="VZU DD BM" number="1">
              <RESULTS>
                <RESULT eventid="1140" reactiontime="+93" status="EXH" swimtime="00:05:24.16" resultid="29383" entrytime="00:05:19.66">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.56" />
                    <SPLIT distance="100" swimtime="00:01:20.67" />
                    <SPLIT distance="150" swimtime="00:01:59.47" />
                    <SPLIT distance="200" swimtime="00:02:42.57" />
                    <SPLIT distance="250" swimtime="00:03:23.38" />
                    <SPLIT distance="300" swimtime="00:04:04.97" />
                    <SPLIT distance="350" swimtime="00:04:41.95" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="29316" number="1" reactiontime="+93" />
                    <RELAYPOSITION athleteid="29279" number="2" reactiontime="+21" />
                    <RELAYPOSITION athleteid="29309" number="3" reactiontime="+95" />
                    <RELAYPOSITION athleteid="29273" number="4" reactiontime="-3" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="13" agetotalmin="12" gender="F" name="VZU DD" number="2">
              <RESULTS>
                <RESULT comment="E1 - Te vroeg overgenomen, waarna niet teruggekeerd naar de bassinwand om opnieuw te vertrekken, 3e te vroeg overgenomen" eventid="1217" reactiontime="+109" status="DSQ" swimtime="00:05:08.16" resultid="29380" entrytime="00:05:12.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.86" />
                    <SPLIT distance="100" swimtime="00:01:24.94" />
                    <SPLIT distance="150" swimtime="00:01:59.53" />
                    <SPLIT distance="200" swimtime="00:02:39.06" />
                    <SPLIT distance="250" swimtime="00:03:13.97" />
                    <SPLIT distance="300" swimtime="00:03:50.65" />
                    <SPLIT distance="350" swimtime="00:04:29.38" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="29316" number="1" reactiontime="+109" status="DSQ" />
                    <RELAYPOSITION athleteid="29279" number="2" reactiontime="+18" status="DSQ" />
                    <RELAYPOSITION athleteid="29273" number="3" reactiontime="-14" status="DSQ" />
                    <RELAYPOSITION athleteid="29309" number="4" reactiontime="+69" status="DSQ" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="13" agetotalmin="12" gender="F" name="VZU DD" number="2">
              <RESULTS>
                <RESULT eventid="26758" reactiontime="+138" swimtime="00:02:12.17" resultid="29381" entrytime="00:02:10.48">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.77" />
                    <SPLIT distance="100" swimtime="00:01:08.67" />
                    <SPLIT distance="150" swimtime="00:01:42.14" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="29316" number="1" reactiontime="+138" />
                    <RELAYPOSITION athleteid="29279" number="2" reactiontime="+15" />
                    <RELAYPOSITION athleteid="29309" number="3" reactiontime="+78" />
                    <RELAYPOSITION athleteid="29273" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="34" agetotalmin="18" gender="X" name="VZU GA" number="1">
              <RESULTS>
                <RESULT eventid="1210" reactiontime="+97" swimtime="00:01:20.67" resultid="29382" entrytime="00:01:21.22">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:20.30" />
                    <SPLIT distance="100" swimtime="00:00:40.03" />
                    <SPLIT distance="150" swimtime="00:01:01.74" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="29323" number="1" reactiontime="+97" />
                    <RELAYPOSITION athleteid="29328" number="2" />
                    <RELAYPOSITION athleteid="29297" number="3" />
                    <RELAYPOSITION athleteid="29350" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="34" agemin="18" agetotalmax="-1" agetotalmin="-1" gender="X" name="VZU GA" number="2">
              <RESULTS>
                <RESULT eventid="1140" reactiontime="+92" swimtime="00:03:52.15" resultid="29384" entrytime="00:03:45.17">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.58" />
                    <SPLIT distance="100" swimtime="00:01:01.32" />
                    <SPLIT distance="150" swimtime="00:01:28.56" />
                    <SPLIT distance="200" swimtime="00:01:58.15" />
                    <SPLIT distance="250" swimtime="00:02:26.04" />
                    <SPLIT distance="300" swimtime="00:02:57.59" />
                    <SPLIT distance="350" swimtime="00:03:23.64" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="29342" number="1" reactiontime="+92" />
                    <RELAYPOSITION athleteid="29328" number="2" reactiontime="+25" />
                    <RELAYPOSITION athleteid="29362" number="3" reactiontime="+37" />
                    <RELAYPOSITION athleteid="29350" number="4" reactiontime="+17" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="34" agemin="18" agetotalmax="-1" agetotalmin="-1" gender="X" name="VZU GA BM" number="3">
              <RESULTS>
                <RESULT comment="A3 - De aangegeven zwemwijze niet uitgevoerd (oa duiken)" eventid="1140" reactiontime="+96" status="DSQ" swimtime="00:04:44.51" resultid="29385" entrytime="00:04:48.15">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.03" />
                    <SPLIT distance="100" swimtime="00:01:08.42" />
                    <SPLIT distance="150" swimtime="00:01:36.90" />
                    <SPLIT distance="200" swimtime="00:02:12.77" />
                    <SPLIT distance="250" swimtime="00:02:52.93" />
                    <SPLIT distance="300" swimtime="00:03:40.50" />
                    <SPLIT distance="350" swimtime="00:04:10.36" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="29302" number="1" reactiontime="+96" status="DSQ" />
                    <RELAYPOSITION athleteid="29335" number="2" reactiontime="+55" status="DSQ" />
                    <RELAYPOSITION athleteid="29359" number="3" reactiontime="+50" status="DSQ" />
                    <RELAYPOSITION athleteid="29297" number="4" reactiontime="+26" status="DSQ" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
          <OFFICIALS>
            <OFFICIAL officialid="2148" firstname="Edwin" grade="Tijdwaarnemer" lastname="Neehus" nation="NED" />
            <OFFICIAL officialid="21300" firstname="Femma" gender="F" grade="Organisatie" lastname="Neehus" nation="NED" />
            <OFFICIAL officialid="21331" firstname="Andine" gender="F" grade="voorstart" lastname="Haazebroek" nation="NED" />
            <OFFICIAL officialid="28781" firstname="Mirjam" gender="F" grade="Medailles" lastname="Jansen" nation="NED" />
            <OFFICIAL officialid="2147" firstname="Dick" gender="M" grade="Starter" lastname="Kuin" nation="NED" />
            <OFFICIAL officialid="3073" firstname="Ande" gender="F" grade="Ploegleider" lastname="Raadschelders" nameprefix=" " nation="NED" />
            <OFFICIAL officialid="23068" firstname="Ytje" gender="F" grade="Lijnrechter" lastname="Munke" nation="NED" />
            <OFFICIAL officialid="5128" firstname="Peter" grade="Tijdwaarnemer" lastname="Raadschelders" nation="NED" />
            <OFFICIAL officialid="28808" firstname="Friso" gender="M" grade="Ploegleider" lastname="Zandwijk" nation="NED" />
            <OFFICIAL officialid="4863" firstname="Jessica" gender="F" grade="Tijdwaarnemer" lastname="Bohm" nation="NED" />
            <OFFICIAL officialid="2149" firstname="Karin" gender="F" grade="Directeur NK" lastname="Neehus" nation="NED" />
          </OFFICIALS>
        </CLUB>
        <CLUB type="CLUB" clubid="28819" name="MET INSCHRIJVINGEN" shortname="MET ">
          <OFFICIALS>
            <OFFICIAL officialid="28821" firstname="BUITENLANDSE " gender="M" grade="MET INSCHRIJVINGEN" lastname="TEAMS" />
            <OFFICIAL officialid="28818" firstname="Nederlandse " gender="M" grade="MET INSCHRIJVINGEN" lastname="Teams" />
          </OFFICIALS>
        </CLUB>
        <CLUB type="CLUB" code="RBT98" nation="NED" clubid="18969" name="Rbt &apos;98">
          <COACHES>
            <COACH firstname="Ferry" gender="M" lastname="Hoogedoorn" nation="NED" type="STAFF" />
          </COACHES>
          <OFFICIALS>
            <OFFICIAL officialid="27733" firstname="Ferry" gender="M" grade="Ploegleider" lastname="Hoogedoorn" nation="NED" />
          </OFFICIALS>
        </CLUB>
        <CLUB type="CLUB" code="FREIBURG" nation="GER" clubid="26906" name="SSV Freiburg">
          <OFFICIALS>
            <OFFICIAL officialid="27691" firstname="Sascha" gender="M" grade="Team Captain" lastname="Schmidt" nation="GER" />
          </OFFICIALS>
        </CLUB>
        <CLUB type="CLUB" code="BTSC" nation="GER" clubid="27600" name="Binger Tauchsportclub eV" shortname="Binger TSC">
          <ATHLETES>
            <ATHLETE firstname="Ben" lastname="Del Sordo" birthdate="2012-01-01" gender="M" nation="GER" license="090191 000612" athleteid="29084">
              <RESULTS>
                <RESULT eventid="1079" points="891" reactiontime="+105" swimtime="00:00:28.85" resultid="29100" entrytime="00:00:30.48" />
                <RESULT eventid="7264" points="604" reactiontime="+108" swimtime="00:06:12.03" resultid="29101" entrytime="00:05:46.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.61" />
                    <SPLIT distance="100" swimtime="00:01:25.92" />
                    <SPLIT distance="150" swimtime="00:02:14.05" />
                    <SPLIT distance="200" swimtime="00:03:05.36" />
                    <SPLIT distance="250" swimtime="00:03:57.60" />
                    <SPLIT distance="300" swimtime="00:04:50.03" />
                    <SPLIT distance="350" swimtime="00:05:35.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="7295" points="830" reactiontime="+107" swimtime="00:01:08.94" resultid="29102" entrytime="00:01:09.84">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="24862" points="631" reactiontime="+100" swimtime="00:02:41.02" resultid="29103" entrytime="00:02:38.13">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.36" />
                    <SPLIT distance="100" swimtime="00:01:20.63" />
                    <SPLIT distance="150" swimtime="00:02:05.95" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Paul" lastname="Funke" birthdate="2008-01-01" gender="M" nation="GER" license="090191 000575" athleteid="29086">
              <RESULTS>
                <RESULT eventid="1079" points="687" reactiontime="+110" swimtime="00:00:23.47" resultid="29110" entrytime="00:00:22.87" />
                <RESULT eventid="7264" points="741" reactiontime="+118" swimtime="00:04:20.13" resultid="29112" entrytime="00:04:05.70">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.90" />
                    <SPLIT distance="100" swimtime="00:00:58.31" />
                    <SPLIT distance="150" swimtime="00:01:31.24" />
                    <SPLIT distance="200" swimtime="00:02:05.05" />
                    <SPLIT distance="250" swimtime="00:02:39.83" />
                    <SPLIT distance="300" swimtime="00:03:14.63" />
                    <SPLIT distance="350" swimtime="00:03:48.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1153" status="WDR" swimtime="00:00:00.00" resultid="29113" entrytime="00:00:24.42" />
                <RESULT eventid="16574" points="900" reactiontime="+112" swimtime="00:08:58.96" resultid="29114" entrytime="00:08:41.97">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.17" />
                    <SPLIT distance="100" swimtime="00:01:00.35" />
                    <SPLIT distance="150" swimtime="00:01:33.74" />
                    <SPLIT distance="200" swimtime="00:02:07.43" />
                    <SPLIT distance="250" swimtime="00:02:41.60" />
                    <SPLIT distance="300" swimtime="00:03:16.02" />
                    <SPLIT distance="350" swimtime="00:03:50.38" />
                    <SPLIT distance="400" swimtime="00:04:24.87" />
                    <SPLIT distance="450" swimtime="00:04:59.51" />
                    <SPLIT distance="500" swimtime="00:05:34.14" />
                    <SPLIT distance="550" swimtime="00:06:08.73" />
                    <SPLIT distance="600" swimtime="00:06:43.85" />
                    <SPLIT distance="650" swimtime="00:07:18.29" />
                    <SPLIT distance="700" swimtime="00:07:53.01" />
                    <SPLIT distance="750" swimtime="00:08:26.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="7295" points="689" reactiontime="+105" swimtime="00:00:51.43" resultid="29115" entrytime="00:00:51.03">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:24.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="24862" points="702" reactiontime="+104" swimtime="00:01:58.90" resultid="29116" entrytime="00:01:54.16">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.00" />
                    <SPLIT distance="100" swimtime="00:00:56.35" />
                    <SPLIT distance="150" swimtime="00:01:27.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="18215" points="729" reactiontime="+100" swimtime="00:17:42.87" resultid="29468" entrytime="00:17:16.08">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.02" />
                    <SPLIT distance="100" swimtime="00:01:03.88" />
                    <SPLIT distance="150" swimtime="00:01:39.83" />
                    <SPLIT distance="200" swimtime="00:02:16.22" />
                    <SPLIT distance="250" swimtime="00:02:52.55" />
                    <SPLIT distance="300" swimtime="00:03:28.44" />
                    <SPLIT distance="350" swimtime="00:04:05.53" />
                    <SPLIT distance="400" swimtime="00:04:41.87" />
                    <SPLIT distance="450" swimtime="00:05:18.09" />
                    <SPLIT distance="500" swimtime="00:05:53.78" />
                    <SPLIT distance="550" swimtime="00:06:29.26" />
                    <SPLIT distance="600" swimtime="00:07:05.22" />
                    <SPLIT distance="650" swimtime="00:07:40.67" />
                    <SPLIT distance="700" swimtime="00:08:16.09" />
                    <SPLIT distance="750" swimtime="00:08:50.95" />
                    <SPLIT distance="800" swimtime="00:09:26.20" />
                    <SPLIT distance="850" swimtime="00:10:02.31" />
                    <SPLIT distance="900" swimtime="00:10:37.78" />
                    <SPLIT distance="950" swimtime="00:11:13.37" />
                    <SPLIT distance="1000" swimtime="00:11:49.43" />
                    <SPLIT distance="1050" swimtime="00:12:25.35" />
                    <SPLIT distance="1100" swimtime="00:13:01.33" />
                    <SPLIT distance="1150" swimtime="00:13:37.58" />
                    <SPLIT distance="1200" swimtime="00:14:13.60" />
                    <SPLIT distance="1250" swimtime="00:14:48.63" />
                    <SPLIT distance="1300" swimtime="00:15:24.48" />
                    <SPLIT distance="1350" swimtime="00:16:00.88" />
                    <SPLIT distance="1400" swimtime="00:16:37.44" />
                    <SPLIT distance="1450" swimtime="00:17:09.57" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Florian" lastname="Funke" birthdate="2010-01-01" gender="M" nation="GER" license="090191 000574" athleteid="29087">
              <RESULTS>
                <RESULT eventid="1079" points="712" reactiontime="+89" swimtime="00:00:26.39" resultid="29117" entrytime="00:00:25.51" />
                <RESULT eventid="7264" points="822" reactiontime="+104" swimtime="00:04:49.89" resultid="29119" entrytime="00:04:29.91">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.08" />
                    <SPLIT distance="100" swimtime="00:01:08.29" />
                    <SPLIT distance="150" swimtime="00:01:45.68" />
                    <SPLIT distance="200" swimtime="00:02:23.89" />
                    <SPLIT distance="250" swimtime="00:03:02.90" />
                    <SPLIT distance="300" swimtime="00:03:38.68" />
                    <SPLIT distance="350" swimtime="00:04:14.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="16574" points="742" reactiontime="+111" swimtime="00:10:08.18" resultid="29120" entrytime="00:09:47.40">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.38" />
                    <SPLIT distance="100" swimtime="00:01:11.07" />
                    <SPLIT distance="150" swimtime="00:01:49.66" />
                    <SPLIT distance="200" swimtime="00:02:29.42" />
                    <SPLIT distance="250" swimtime="00:03:09.09" />
                    <SPLIT distance="300" swimtime="00:03:48.38" />
                    <SPLIT distance="350" swimtime="00:04:28.42" />
                    <SPLIT distance="400" swimtime="00:05:06.18" />
                    <SPLIT distance="450" swimtime="00:05:43.81" />
                    <SPLIT distance="500" swimtime="00:06:21.63" />
                    <SPLIT distance="550" swimtime="00:06:59.03" />
                    <SPLIT distance="600" swimtime="00:07:37.65" />
                    <SPLIT distance="650" swimtime="00:08:17.38" />
                    <SPLIT distance="700" swimtime="00:08:55.54" />
                    <SPLIT distance="750" swimtime="00:09:33.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="7295" points="688" reactiontime="+89" swimtime="00:01:01.67" resultid="29121" entrytime="00:00:58.07">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="18215" reactiontime="+117" swimtime="00:20:07.40" resultid="29467" entrytime="00:21:00.74">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.18" />
                    <SPLIT distance="100" swimtime="00:01:16.09" />
                    <SPLIT distance="150" swimtime="00:01:55.92" />
                    <SPLIT distance="200" swimtime="00:02:35.05" />
                    <SPLIT distance="250" swimtime="00:03:14.70" />
                    <SPLIT distance="300" swimtime="00:03:54.27" />
                    <SPLIT distance="350" swimtime="00:04:35.63" />
                    <SPLIT distance="400" swimtime="00:05:18.77" />
                    <SPLIT distance="450" swimtime="00:06:01.69" />
                    <SPLIT distance="500" swimtime="00:06:44.50" />
                    <SPLIT distance="550" swimtime="00:07:28.88" />
                    <SPLIT distance="600" swimtime="00:08:08.79" />
                    <SPLIT distance="650" swimtime="00:08:52.36" />
                    <SPLIT distance="700" swimtime="00:09:35.19" />
                    <SPLIT distance="750" swimtime="00:10:17.59" />
                    <SPLIT distance="800" swimtime="00:10:59.74" />
                    <SPLIT distance="850" swimtime="00:11:42.33" />
                    <SPLIT distance="900" swimtime="00:12:26.83" />
                    <SPLIT distance="950" swimtime="00:13:05.88" />
                    <SPLIT distance="1000" swimtime="00:13:45.79" />
                    <SPLIT distance="1050" swimtime="00:14:24.76" />
                    <SPLIT distance="1100" swimtime="00:15:04.66" />
                    <SPLIT distance="1150" swimtime="00:15:43.90" />
                    <SPLIT distance="1200" swimtime="00:16:22.31" />
                    <SPLIT distance="1250" swimtime="00:17:01.38" />
                    <SPLIT distance="1300" swimtime="00:17:40.45" />
                    <SPLIT distance="1350" swimtime="00:18:20.97" />
                    <SPLIT distance="1400" swimtime="00:18:56.12" />
                    <SPLIT distance="1450" swimtime="00:19:33.87" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Stella" lastname="Jöckel" birthdate="2007-01-01" gender="F" nation="GER" license="090191 000586" athleteid="29083">
              <RESULTS>
                <RESULT eventid="1053" points="290" reactiontime="+102" swimtime="00:00:31.12" resultid="29094" entrytime="00:00:32.72" />
                <RESULT eventid="7278" points="303" reactiontime="+98" swimtime="00:05:36.01" resultid="29095" entrytime="00:05:57.01">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.85" />
                    <SPLIT distance="100" swimtime="00:01:16.96" />
                    <SPLIT distance="150" swimtime="00:02:00.81" />
                    <SPLIT distance="200" swimtime="00:02:46.03" />
                    <SPLIT distance="250" swimtime="00:03:30.09" />
                    <SPLIT distance="300" swimtime="00:04:15.21" />
                    <SPLIT distance="350" swimtime="00:04:58.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1147" points="246" reactiontime="+95" swimtime="00:00:30.61" resultid="29096" entrytime="00:00:33.64" />
                <RESULT eventid="1158" points="268" reactiontime="+103" swimtime="00:12:05.52" resultid="29097" entrytime="00:12:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.01" />
                    <SPLIT distance="100" swimtime="00:01:23.58" />
                    <SPLIT distance="150" swimtime="00:02:10.20" />
                    <SPLIT distance="200" swimtime="00:02:56.08" />
                    <SPLIT distance="250" swimtime="00:03:42.52" />
                    <SPLIT distance="300" swimtime="00:04:28.86" />
                    <SPLIT distance="350" swimtime="00:05:15.89" />
                    <SPLIT distance="400" swimtime="00:06:04.47" />
                    <SPLIT distance="450" swimtime="00:06:52.23" />
                    <SPLIT distance="500" swimtime="00:07:41.36" />
                    <SPLIT distance="550" swimtime="00:08:30.40" />
                    <SPLIT distance="600" swimtime="00:09:17.70" />
                    <SPLIT distance="650" swimtime="00:10:03.85" />
                    <SPLIT distance="700" swimtime="00:10:48.90" />
                    <SPLIT distance="750" swimtime="00:11:28.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="7287" points="220" reactiontime="+106" swimtime="00:01:16.60" resultid="29098" entrytime="00:01:11.39">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="24851" status="WDR" swimtime="00:00:00.00" resultid="29099" entrytime="00:02:47.49" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lisa" lastname="Walter" birthdate="1997-08-29" gender="F" nation="GER" license="090191 000278" athleteid="27601">
              <RESULTS>
                <RESULT eventid="1053" points="458" reactiontime="+91" swimtime="00:00:25.89" resultid="29091" entrytime="00:00:24.97" />
                <RESULT eventid="1093" points="416" reactiontime="+108" swimtime="00:20:10.70" resultid="29092" entrytime="00:19:19.22">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.35" />
                    <SPLIT distance="100" swimtime="00:01:13.06" />
                    <SPLIT distance="150" swimtime="00:01:52.26" />
                    <SPLIT distance="200" swimtime="00:02:32.48" />
                    <SPLIT distance="250" swimtime="00:03:12.60" />
                    <SPLIT distance="300" swimtime="00:03:53.10" />
                    <SPLIT distance="350" swimtime="00:04:32.83" />
                    <SPLIT distance="400" swimtime="00:05:12.79" />
                    <SPLIT distance="450" swimtime="00:05:53.98" />
                    <SPLIT distance="500" swimtime="00:06:34.67" />
                    <SPLIT distance="550" swimtime="00:07:16.25" />
                    <SPLIT distance="600" swimtime="00:07:56.57" />
                    <SPLIT distance="650" swimtime="00:08:38.28" />
                    <SPLIT distance="700" swimtime="00:09:19.05" />
                    <SPLIT distance="750" swimtime="00:10:00.66" />
                    <SPLIT distance="800" swimtime="00:10:42.01" />
                    <SPLIT distance="850" swimtime="00:11:23.27" />
                    <SPLIT distance="900" swimtime="00:12:04.66" />
                    <SPLIT distance="950" swimtime="00:12:46.21" />
                    <SPLIT distance="1000" swimtime="00:13:27.32" />
                    <SPLIT distance="1050" swimtime="00:14:08.92" />
                    <SPLIT distance="1100" swimtime="00:14:50.63" />
                    <SPLIT distance="1150" swimtime="00:15:32.32" />
                    <SPLIT distance="1200" swimtime="00:16:13.28" />
                    <SPLIT distance="1250" swimtime="00:16:52.94" />
                    <SPLIT distance="1300" swimtime="00:17:33.36" />
                    <SPLIT distance="1350" swimtime="00:18:14.76" />
                    <SPLIT distance="1400" swimtime="00:18:54.78" />
                    <SPLIT distance="1450" swimtime="00:19:32.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="7278" points="571" reactiontime="+103" swimtime="00:04:30.14" resultid="29093" entrytime="00:04:16.96">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.90" />
                    <SPLIT distance="100" swimtime="00:01:01.86" />
                    <SPLIT distance="150" swimtime="00:01:36.96" />
                    <SPLIT distance="200" swimtime="00:02:12.24" />
                    <SPLIT distance="250" swimtime="00:02:47.06" />
                    <SPLIT distance="300" swimtime="00:03:21.85" />
                    <SPLIT distance="350" swimtime="00:03:56.52" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Julia" lastname="Walter" birthdate="2004-01-01" gender="F" nation="GER" license="090191 000278" athleteid="29082">
              <RESULTS>
                <RESULT eventid="1053" points="544" reactiontime="+95" swimtime="00:00:24.45" resultid="29088" entrytime="00:00:22.95" />
                <RESULT eventid="1093" points="340" reactiontime="+87" swimtime="00:21:34.18" resultid="29089" entrytime="00:21:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.26" />
                    <SPLIT distance="100" swimtime="00:01:14.69" />
                    <SPLIT distance="150" swimtime="00:01:57.19" />
                    <SPLIT distance="200" swimtime="00:02:40.18" />
                    <SPLIT distance="250" swimtime="00:03:19.27" />
                    <SPLIT distance="300" swimtime="00:04:04.88" />
                    <SPLIT distance="350" swimtime="00:04:49.27" />
                    <SPLIT distance="400" swimtime="00:05:35.93" />
                    <SPLIT distance="450" swimtime="00:06:21.44" />
                    <SPLIT distance="500" swimtime="00:07:03.36" />
                    <SPLIT distance="550" swimtime="00:07:49.88" />
                    <SPLIT distance="600" swimtime="00:08:36.60" />
                    <SPLIT distance="650" swimtime="00:09:22.35" />
                    <SPLIT distance="700" swimtime="00:10:08.27" />
                    <SPLIT distance="750" swimtime="00:10:54.53" />
                    <SPLIT distance="800" swimtime="00:11:40.95" />
                    <SPLIT distance="850" swimtime="00:12:28.47" />
                    <SPLIT distance="900" swimtime="00:13:15.75" />
                    <SPLIT distance="950" swimtime="00:14:02.65" />
                    <SPLIT distance="1000" swimtime="00:14:44.63" />
                    <SPLIT distance="1050" swimtime="00:15:30.64" />
                    <SPLIT distance="1100" swimtime="00:16:14.86" />
                    <SPLIT distance="1150" swimtime="00:16:57.70" />
                    <SPLIT distance="1200" swimtime="00:17:35.80" />
                    <SPLIT distance="1250" swimtime="00:18:19.80" />
                    <SPLIT distance="1300" swimtime="00:19:02.40" />
                    <SPLIT distance="1350" swimtime="00:19:37.68" />
                    <SPLIT distance="1400" swimtime="00:20:19.79" />
                    <SPLIT distance="1450" swimtime="00:20:55.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="7278" points="644" reactiontime="+101" swimtime="00:04:19.51" resultid="29090" entrytime="00:04:04.35">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.52" />
                    <SPLIT distance="100" swimtime="00:00:57.93" />
                    <SPLIT distance="150" swimtime="00:01:30.28" />
                    <SPLIT distance="200" swimtime="00:02:04.27" />
                    <SPLIT distance="250" swimtime="00:02:38.96" />
                    <SPLIT distance="300" swimtime="00:03:12.86" />
                    <SPLIT distance="350" swimtime="00:03:46.64" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jan" lastname="Blaszczyk" birthdate="2006-01-01" gender="M" nation="GER" license="090191 000554" athleteid="29085">
              <RESULTS>
                <RESULT eventid="1079" points="756" reactiontime="+133" swimtime="00:00:20.57" resultid="29104" entrytime="00:00:21.94" />
                <RESULT eventid="7264" points="590" reactiontime="+92" swimtime="00:04:10.31" resultid="29105" entrytime="00:04:07.09">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:24.76" />
                    <SPLIT distance="100" swimtime="00:00:53.20" />
                    <SPLIT distance="150" swimtime="00:01:24.17" />
                    <SPLIT distance="200" swimtime="00:01:56.93" />
                    <SPLIT distance="250" swimtime="00:02:30.52" />
                    <SPLIT distance="300" swimtime="00:03:03.93" />
                    <SPLIT distance="350" swimtime="00:03:37.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1153" points="679" reactiontime="+108" swimtime="00:00:19.28" resultid="29106" entrytime="00:00:20.01" />
                <RESULT eventid="16574" points="623" reactiontime="+101" swimtime="00:08:41.53" resultid="29107" entrytime="00:08:47.09">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.52" />
                    <SPLIT distance="100" swimtime="00:00:56.56" />
                    <SPLIT distance="150" swimtime="00:01:28.03" />
                    <SPLIT distance="200" swimtime="00:02:00.01" />
                    <SPLIT distance="250" swimtime="00:02:32.61" />
                    <SPLIT distance="300" swimtime="00:03:05.47" />
                    <SPLIT distance="350" swimtime="00:03:39.28" />
                    <SPLIT distance="400" swimtime="00:04:13.28" />
                    <SPLIT distance="450" swimtime="00:04:47.89" />
                    <SPLIT distance="500" swimtime="00:05:21.74" />
                    <SPLIT distance="550" swimtime="00:05:55.77" />
                    <SPLIT distance="600" swimtime="00:06:29.52" />
                    <SPLIT distance="650" swimtime="00:07:03.91" />
                    <SPLIT distance="700" swimtime="00:07:37.62" />
                    <SPLIT distance="750" swimtime="00:08:10.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="7295" points="667" reactiontime="+106" swimtime="00:00:46.71" resultid="29108" entrytime="00:00:49.48">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:21.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="24862" points="774" reactiontime="+106" swimtime="00:01:51.67" resultid="29109" entrytime="00:01:54.78">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.35" />
                    <SPLIT distance="100" swimtime="00:00:53.98" />
                    <SPLIT distance="150" swimtime="00:01:23.52" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="17" agetotalmin="16" gender="M" name="Binger TC HB" number="1">
              <RESULTS>
                <RESULT comment="B2 - Na start- en/of keerpunt meer dan 15 meter onder water gezwommen" eventid="26768" reactiontime="+98" status="DSQ" swimtime="00:01:39.06" resultid="29122" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:20.57" />
                    <SPLIT distance="100" swimtime="00:00:46.92" />
                    <SPLIT distance="150" swimtime="00:01:09.92" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="29085" number="1" reactiontime="+98" status="DSQ" />
                    <RELAYPOSITION athleteid="29087" number="2" reactiontime="+64" status="DSQ" />
                    <RELAYPOSITION athleteid="29086" number="3" reactiontime="+54" status="DSQ" />
                    <RELAYPOSITION athleteid="29084" number="4" reactiontime="+81" status="DSQ" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="17" agetotalmin="16" gender="M" name="Binger TC HB" number="1">
              <RESULTS>
                <RESULT eventid="24873" reactiontime="+101" swimtime="00:03:49.67" resultid="29123" entrytime="00:03:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:22.07" />
                    <SPLIT distance="100" swimtime="00:00:46.46" />
                    <SPLIT distance="150" swimtime="00:01:13.81" />
                    <SPLIT distance="200" swimtime="00:01:46.27" />
                    <SPLIT distance="250" swimtime="00:02:10.71" />
                    <SPLIT distance="300" swimtime="00:02:39.11" />
                    <SPLIT distance="350" swimtime="00:03:12.66" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="29085" number="1" reactiontime="+101" />
                    <RELAYPOSITION athleteid="29087" number="2" reactiontime="+56" />
                    <RELAYPOSITION athleteid="29086" number="3" reactiontime="+69" />
                    <RELAYPOSITION athleteid="29084" number="4" reactiontime="+77" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
          <OFFICIALS>
            <OFFICIAL officialid="27683" firstname="Sandra" gender="F" grade="Team Captain" lastname="Funcke" nation="GER" />
          </OFFICIALS>
        </CLUB>
        <CLUB type="CLUB" code="TSCR1957" nation="GER" clubid="22578" name="TSC Rostock 1957" />
        <CLUB type="CLUB" code="CPB RENNES" nation="FRA" clubid="27825" name="Cercle Paul Bert Rennes" shortname="CPB Rennes">
          <ATHLETES>
            <ATHLETE firstname="Anais" lastname="Verger" birthdate="2000-01-01" gender="F" nation="FRA" license="A-18-797507" athleteid="28936">
              <RESULTS>
                <RESULT comment="backup tijd" eventid="1053" points="1316" reactiontime="+88" swimtime="00:00:18.21" resultid="28937" entrytime="00:00:18.93" />
                <RESULT eventid="1120" points="1042" reactiontime="+83" swimtime="00:00:23.01" resultid="28938" entrytime="00:00:22.98" />
                <RESULT comment="Backup tijd" eventid="1147" points="1363" reactiontime="+87" swimtime="00:00:17.00" resultid="28939" entrytime="00:00:17.27" />
                <RESULT eventid="7287" points="1459" reactiontime="+93" swimtime="00:00:40.48" resultid="28940" entrytime="00:00:40.57">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:19.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="24851" points="1328" reactiontime="+92" swimtime="00:01:32.14" resultid="28941" entrytime="00:01:31.66">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:21.71" />
                    <SPLIT distance="100" swimtime="00:00:44.60" />
                    <SPLIT distance="150" swimtime="00:01:08.54" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <OFFICIALS>
            <OFFICIAL officialid="27826" firstname="Hugues" gender="M" grade="Team Captain" lastname="Brilhault" nation="FRA" />
          </OFFICIALS>
        </CLUB>
        <CLUB type="CLUB" nation="NED" clubid="22896" name="Unattached">
          <OFFICIALS>
            <OFFICIAL officialid="1508" firstname="Lonny" gender="F" grade="Vz. Kamprechter" lastname="Hendriks" nation="NED" />
            <OFFICIAL officialid="1510" firstname="Roland" gender="M" grade="Starter" lastname="Kanters" nation="NED" />
            <OFFICIAL officialid="1547" firstname="Lonny" gender="F" grade=" VK, Kamprechter, Ti" lastname="Hendriks" nation="NED" />
            <OFFICIAL officialid="3067" firstname="Kees" grade="Secretariaat" lastname="Bom" nation="NED" />
          </OFFICIALS>
        </CLUB>
        <CLUB type="CLUB" code="CAAP" nation="FRA" clubid="24487" name="CAAP" />
        <CLUB type="CLUB" code="DJK-VFR" nation="GER" clubid="22537" name="DJK-VfR Mülheim Saarn">
          <ATHLETES>
            <ATHLETE firstname="Luis" lastname="Grinten" birthdate="2012-08-26" gender="M" nameprefix="van der" nation="GER" license=".80060000533" athleteid="28158">
              <RESULTS>
                <RESULT eventid="1079" points="769" reactiontime="+83" swimtime="00:00:30.31" resultid="28159" entrytime="00:00:32.58" />
                <RESULT eventid="7271" points="872" reactiontime="+104" swimtime="00:02:38.01" resultid="28160" entrytime="00:03:14.25">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.55" />
                    <SPLIT distance="100" swimtime="00:01:15.74" />
                    <SPLIT distance="150" swimtime="00:01:59.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1127" points="948" reactiontime="+88" swimtime="00:00:30.63" resultid="28161" entrytime="00:00:33.78" />
                <RESULT eventid="7264" points="760" reactiontime="+115" swimtime="00:05:44.70" resultid="28162" entrytime="00:05:48.87">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.50" />
                    <SPLIT distance="100" swimtime="00:01:18.08" />
                    <SPLIT distance="200" swimtime="00:02:46.28" />
                    <SPLIT distance="250" swimtime="00:03:31.01" />
                    <SPLIT distance="300" swimtime="00:04:16.94" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rebecca" lastname="Howe" birthdate="2009-09-14" gender="F" nation="GER" license=".80060000534" athleteid="28153">
              <RESULTS>
                <RESULT eventid="1053" points="440" reactiontime="+145" swimtime="00:00:28.15" resultid="28154" entrytime="00:00:30.58" />
                <RESULT eventid="7254" points="622" reactiontime="+115" swimtime="00:02:28.44" resultid="28155" entrytime="00:03:02.32">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.57" />
                    <SPLIT distance="100" swimtime="00:01:10.71" />
                    <SPLIT distance="150" swimtime="00:01:51.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1120" points="671" reactiontime="+101" swimtime="00:00:28.36" resultid="28156" entrytime="00:00:31.67" />
                <RESULT eventid="7278" points="294" reactiontime="+133" swimtime="00:05:47.89" resultid="28157" entrytime="00:04:52.06">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.82" />
                    <SPLIT distance="100" swimtime="00:01:15.20" />
                    <SPLIT distance="150" swimtime="00:01:58.97" />
                    <SPLIT distance="200" swimtime="00:02:47.24" />
                    <SPLIT distance="250" swimtime="00:03:32.68" />
                    <SPLIT distance="300" swimtime="00:04:14.80" />
                    <SPLIT distance="350" swimtime="00:05:03.80" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marvin" lastname="Venohr" birthdate="2000-07-17" gender="M" nation="GER" license=".80060000541" athleteid="28163">
              <RESULTS>
                <RESULT eventid="1079" points="443" reactiontime="+109" swimtime="00:00:22.23" resultid="28164" entrytime="00:00:22.98" />
                <RESULT eventid="7271" points="669" reactiontime="+105" swimtime="00:02:04.56" resultid="28165" entrytime="00:02:02.25">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.86" />
                    <SPLIT distance="100" swimtime="00:00:58.37" />
                    <SPLIT distance="150" swimtime="00:01:31.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="7264" points="485" reactiontime="+120" swimtime="00:04:10.06" resultid="28166" entrytime="00:04:09.64">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.54" />
                    <SPLIT distance="100" swimtime="00:00:59.24" />
                    <SPLIT distance="150" swimtime="00:01:31.06" />
                    <SPLIT distance="200" swimtime="00:02:03.67" />
                    <SPLIT distance="250" swimtime="00:02:36.82" />
                    <SPLIT distance="300" swimtime="00:03:09.41" />
                    <SPLIT distance="350" swimtime="00:03:41.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1153" points="447" reactiontime="+110" swimtime="00:00:20.67" resultid="28167" entrytime="00:00:22.23" />
                <RESULT eventid="1175" points="603" reactiontime="+98" swimtime="00:00:54.63" resultid="28168" entrytime="00:00:53.31">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="7295" points="508" reactiontime="+111" swimtime="00:00:49.39" resultid="28169" entrytime="00:00:48.51">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:23.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="24862" points="546" reactiontime="+114" swimtime="00:01:52.42" resultid="28170" entrytime="00:01:55.25">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.58" />
                    <SPLIT distance="100" swimtime="00:00:53.39" />
                    <SPLIT distance="150" swimtime="00:01:23.15" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Phil Jason" lastname="Bieler" birthdate="2005-10-10" gender="M" nation="GER" license=".80060000457" athleteid="28171">
              <RESULTS>
                <RESULT eventid="1079" points="732" reactiontime="+94" swimtime="00:00:18.80" resultid="28172" entrytime="00:00:19.61" />
                <RESULT eventid="26746" points="1017" reactiontime="+110" swimtime="00:06:44.31" resultid="28173" entrytime="00:07:05.41">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:21.51" />
                    <SPLIT distance="100" swimtime="00:00:44.83" />
                    <SPLIT distance="150" swimtime="00:01:09.64" />
                    <SPLIT distance="200" swimtime="00:01:35.11" />
                    <SPLIT distance="250" swimtime="00:02:00.60" />
                    <SPLIT distance="300" swimtime="00:02:27.00" />
                    <SPLIT distance="350" swimtime="00:02:52.86" />
                    <SPLIT distance="400" swimtime="00:03:18.67" />
                    <SPLIT distance="450" swimtime="00:03:44.89" />
                    <SPLIT distance="500" swimtime="00:04:11.33" />
                    <SPLIT distance="550" swimtime="00:04:37.51" />
                    <SPLIT distance="600" swimtime="00:05:03.10" />
                    <SPLIT distance="650" swimtime="00:05:29.04" />
                    <SPLIT distance="700" swimtime="00:05:54.83" />
                    <SPLIT distance="750" swimtime="00:06:20.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1114" points="983" reactiontime="+107" swimtime="00:03:13.92" resultid="28174" entrytime="00:03:12.39">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:21.10" />
                    <SPLIT distance="100" swimtime="00:00:44.20" />
                    <SPLIT distance="150" swimtime="00:01:08.86" />
                    <SPLIT distance="200" swimtime="00:01:34.17" />
                    <SPLIT distance="250" swimtime="00:01:59.52" />
                    <SPLIT distance="300" swimtime="00:02:24.53" />
                    <SPLIT distance="350" swimtime="00:02:50.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="16574" points="917" reactiontime="+91" swimtime="00:07:04.81" resultid="28175" entrytime="00:07:09.11">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:21.88" />
                    <SPLIT distance="100" swimtime="00:00:47.23" />
                    <SPLIT distance="150" swimtime="00:01:14.13" />
                    <SPLIT distance="200" swimtime="00:01:41.24" />
                    <SPLIT distance="250" swimtime="00:02:08.34" />
                    <SPLIT distance="300" swimtime="00:02:35.38" />
                    <SPLIT distance="350" swimtime="00:03:03.06" />
                    <SPLIT distance="400" swimtime="00:03:30.51" />
                    <SPLIT distance="450" swimtime="00:03:58.04" />
                    <SPLIT distance="500" swimtime="00:04:25.41" />
                    <SPLIT distance="550" swimtime="00:04:52.22" />
                    <SPLIT distance="600" swimtime="00:05:19.55" />
                    <SPLIT distance="650" swimtime="00:05:46.90" />
                    <SPLIT distance="700" swimtime="00:06:14.07" />
                    <SPLIT distance="750" swimtime="00:06:40.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="24862" points="972" reactiontime="+89" swimtime="00:01:32.78" resultid="28176" entrytime="00:01:40.55">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:20.82" />
                    <SPLIT distance="100" swimtime="00:00:44.32" />
                    <SPLIT distance="150" swimtime="00:01:09.32" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Valeria" lastname="Lazarenko" birthdate="2010-04-01" gender="F" nation="UKR" license=".80060000540" athleteid="27074">
              <RESULTS>
                <RESULT eventid="1053" points="1091" reactiontime="+96" swimtime="00:00:22.05" resultid="28149" entrytime="00:00:23.16" />
                <RESULT eventid="7278" points="1578" reactiontime="+101" swimtime="00:03:56.95" resultid="28150" entrytime="00:04:05.64">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.12" />
                    <SPLIT distance="100" swimtime="00:00:54.57" />
                    <SPLIT distance="150" swimtime="00:01:24.79" />
                    <SPLIT distance="200" swimtime="00:01:55.58" />
                    <SPLIT distance="250" swimtime="00:02:26.73" />
                    <SPLIT distance="300" swimtime="00:02:57.84" />
                    <SPLIT distance="350" swimtime="00:03:28.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="7287" status="WDR" swimtime="00:00:00.00" resultid="28151" entrytime="00:00:51.66" />
                <RESULT eventid="1182" status="WDR" swimtime="00:00:00.00" resultid="28152" entrytime="00:00:47.15" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="34" agemin="18" agetotalmax="-1" agetotalmin="-1" gender="X" name="DJK-VFR GA" number="1">
              <RESULTS>
                <RESULT eventid="1140" reactiontime="+89" swimtime="00:03:49.78" resultid="28177" entrytime="00:04:35.72" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:24.18" />
                    <SPLIT distance="100" swimtime="00:00:50.56" />
                    <SPLIT distance="150" swimtime="00:01:18.91" />
                    <SPLIT distance="200" swimtime="00:01:49.44" />
                    <SPLIT distance="250" swimtime="00:02:16.36" />
                    <SPLIT distance="300" swimtime="00:02:45.46" />
                    <SPLIT distance="350" swimtime="00:03:16.16" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="28171" number="1" reactiontime="+89" />
                    <RELAYPOSITION athleteid="27074" number="2" reactiontime="+68" />
                    <RELAYPOSITION athleteid="28163" number="3" reactiontime="+73" />
                    <RELAYPOSITION athleteid="28153" number="4" reactiontime="+57" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
          <OFFICIALS>
            <OFFICIAL officialid="24198" firstname="Leo" gender="M" grade="Team Captain" lastname="Runge" nation="GER" />
            <OFFICIAL officialid="28487" firstname="Karina " gender="M" grade="Tijdwaarnemer in opl" lastname="Lazarenko" nation="GER" />
            <OFFICIAL officialid="23071" firstname="Heike" gender="F" grade="Tijdwaarnemer" lastname="Bieler" nation="GER" />
          </OFFICIALS>
        </CLUB>
        <CLUB type="CLUB" code="CSL" nation="FRA" clubid="26042" name="CS Lorientais" shortname="CSL">
          <OFFICIALS>
            <OFFICIAL officialid="28806" firstname="Olivier" gender="M" grade="Team Captain" lastname="Milleville" nation="FRA" />
          </OFFICIALS>
        </CLUB>
        <CLUB type="CLUB" code="PONTOS" nation="NED" clubid="17046" name="OWT Pontos" shortname="PONTOS">
          <ATHLETES>
            <ATHLETE firstname="Silke" lastname="Geest" birthdate="2008-10-16" gender="F" nameprefix="van der" nation="NED" license="9261622" athleteid="28252">
              <RESULTS>
                <RESULT eventid="1053" points="696" reactiontime="+94" swimtime="00:00:24.17" resultid="28253" entrytime="00:00:25.34" entrycourse="LCM" />
                <RESULT eventid="7254" points="708" reactiontime="+103" swimtime="00:02:22.17" resultid="28254">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.23" />
                    <SPLIT distance="100" swimtime="00:01:05.69" />
                    <SPLIT distance="150" swimtime="00:01:44.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1120" points="669" reactiontime="+104" swimtime="00:00:28.39" resultid="28255" entrytime="00:00:28.41" />
                <RESULT eventid="1147" points="512" reactiontime="+99" swimtime="00:00:24.00" resultid="28256" />
                <RESULT eventid="1168" points="749" reactiontime="+100" swimtime="00:01:02.43" resultid="28257" entrytime="00:01:04.07">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="7287" points="634" reactiontime="+109" swimtime="00:00:55.00" resultid="28258" entrytime="00:00:57.06">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="24851" points="593" reactiontime="+98" swimtime="00:02:06.13" resultid="28259" entrytime="00:02:11.89" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.19" />
                    <SPLIT distance="100" swimtime="00:00:57.15" />
                    <SPLIT distance="150" swimtime="00:01:32.00" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Sanne" lastname="Fuchten" birthdate="2009-12-16" gender="F" nation="NED" license="9228724" athleteid="28246">
              <RESULTS>
                <RESULT eventid="1053" points="305" reactiontime="+98" swimtime="00:00:31.79" resultid="28247" entrytime="00:00:32.67" entrycourse="LCM" />
                <RESULT eventid="7254" points="573" reactiontime="+98" swimtime="00:02:32.54" resultid="28248" entrytime="00:02:46.99" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.49" />
                    <SPLIT distance="100" swimtime="00:01:11.60" />
                    <SPLIT distance="150" swimtime="00:01:52.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1120" points="458" reactiontime="+108" swimtime="00:00:32.19" resultid="28249" entrytime="00:00:32.43" entrycourse="LCM" />
                <RESULT eventid="1168" points="493" reactiontime="+109" swimtime="00:01:11.74" resultid="28250" entrytime="00:01:11.60" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1196" points="683" reactiontime="+115" swimtime="00:05:22.70" resultid="28251" entrytime="00:05:38.13" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.20" />
                    <SPLIT distance="100" swimtime="00:01:18.96" />
                    <SPLIT distance="150" swimtime="00:02:00.10" />
                    <SPLIT distance="200" swimtime="00:02:41.24" />
                    <SPLIT distance="250" swimtime="00:03:22.34" />
                    <SPLIT distance="300" swimtime="00:04:04.05" />
                    <SPLIT distance="350" swimtime="00:04:44.91" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Janneke" lastname="Mandigers" birthdate="2001-04-17" gender="F" nation="NED" license="9013717" athleteid="28282">
              <RESULTS>
                <RESULT eventid="1053" points="518" reactiontime="+107" swimtime="00:00:24.84" resultid="28283" entrytime="00:00:26.40" entrycourse="LCM" />
                <RESULT eventid="7254" points="547" reactiontime="+97" swimtime="00:02:15.09" resultid="28284" entrytime="00:02:21.94" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.78" />
                    <SPLIT distance="100" swimtime="00:01:04.84" />
                    <SPLIT distance="150" swimtime="00:01:40.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1120" points="546" reactiontime="+97" swimtime="00:00:28.54" resultid="28285" entrytime="00:00:29.46" entrycourse="LCM" />
                <RESULT eventid="7278" points="563" reactiontime="+102" swimtime="00:04:31.42" resultid="28286" entrytime="00:04:31.46" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.29" />
                    <SPLIT distance="100" swimtime="00:01:01.82" />
                    <SPLIT distance="150" swimtime="00:01:36.12" />
                    <SPLIT distance="200" swimtime="00:02:11.50" />
                    <SPLIT distance="250" swimtime="00:02:46.52" />
                    <SPLIT distance="300" swimtime="00:03:22.29" />
                    <SPLIT distance="350" swimtime="00:03:58.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1147" points="551" reactiontime="+96" swimtime="00:00:22.98" resultid="28287" entrytime="00:00:24.90" entrycourse="LCM" />
                <RESULT eventid="1158" points="494" reactiontime="+104" swimtime="00:09:52.10" resultid="28288" entrytime="00:09:48.31" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.59" />
                    <SPLIT distance="100" swimtime="00:01:06.53" />
                    <SPLIT distance="150" swimtime="00:01:43.11" />
                    <SPLIT distance="200" swimtime="00:02:20.06" />
                    <SPLIT distance="250" swimtime="00:02:57.60" />
                    <SPLIT distance="300" swimtime="00:03:35.62" />
                    <SPLIT distance="350" swimtime="00:04:13.14" />
                    <SPLIT distance="400" swimtime="00:04:51.20" />
                    <SPLIT distance="450" swimtime="00:05:28.38" />
                    <SPLIT distance="500" swimtime="00:06:05.64" />
                    <SPLIT distance="550" swimtime="00:06:44.11" />
                    <SPLIT distance="600" swimtime="00:07:22.10" />
                    <SPLIT distance="650" swimtime="00:08:00.31" />
                    <SPLIT distance="700" swimtime="00:08:37.71" />
                    <SPLIT distance="750" swimtime="00:09:16.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="7287" points="571" reactiontime="+94" swimtime="00:00:55.35" resultid="28289" entrytime="00:00:59.95" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="24851" points="566" reactiontime="+91" swimtime="00:02:02.41" resultid="28290" entrytime="00:02:07.08" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.31" />
                    <SPLIT distance="100" swimtime="00:00:57.77" />
                    <SPLIT distance="150" swimtime="00:01:30.49" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pien" lastname="Loeffen" birthdate="2010-05-09" gender="F" nation="NED" license="9256869" athleteid="28271">
              <RESULTS>
                <RESULT eventid="1053" points="503" reactiontime="+96" swimtime="00:00:28.53" resultid="28272" entrytime="00:00:29.55" entrycourse="LCM" />
                <RESULT eventid="7254" points="817" reactiontime="+72" swimtime="00:02:24.59" resultid="28273" entrytime="00:02:34.42" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.57" />
                    <SPLIT distance="100" swimtime="00:01:07.43" />
                    <SPLIT distance="150" swimtime="00:01:47.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1120" points="793" reactiontime="+100" swimtime="00:00:29.49" resultid="28274" entrytime="00:00:29.52" entrycourse="LCM" />
                <RESULT eventid="1168" points="713" reactiontime="+100" swimtime="00:01:06.18" resultid="28275" entrytime="00:01:08.06" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1196" points="822" reactiontime="+99" swimtime="00:05:14.72" resultid="28276" entrytime="00:05:37.18" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.96" />
                    <SPLIT distance="100" swimtime="00:01:12.66" />
                    <SPLIT distance="150" swimtime="00:01:52.96" />
                    <SPLIT distance="200" swimtime="00:02:33.96" />
                    <SPLIT distance="250" swimtime="00:03:15.64" />
                    <SPLIT distance="300" swimtime="00:03:57.69" />
                    <SPLIT distance="350" swimtime="00:04:38.60" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Babet" lastname="Fleuren" birthdate="2012-12-22" gender="F" nation="NED" license="9261730" athleteid="28239">
              <RESULTS>
                <RESULT eventid="1053" points="445" reactiontime="+171" swimtime="00:00:33.63" resultid="28240" entrytime="00:00:36.92" entrycourse="LCM" />
                <RESULT eventid="7254" points="589" reactiontime="+112" swimtime="00:03:07.42" resultid="28241" entrytime="00:03:10.93" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.78" />
                    <SPLIT distance="100" swimtime="00:01:26.79" />
                    <SPLIT distance="150" swimtime="00:02:17.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1120" points="570" reactiontime="+115" swimtime="00:00:36.03" resultid="28242" entrytime="00:00:36.80" entrycourse="LCM" />
                <RESULT eventid="1168" points="458" reactiontime="+121" swimtime="00:01:23.66" resultid="28243" entrytime="00:01:26.57" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1196" points="650" reactiontime="+125" swimtime="00:06:29.65" resultid="28244">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.23" />
                    <SPLIT distance="100" swimtime="00:01:25.76" />
                    <SPLIT distance="150" swimtime="00:02:14.96" />
                    <SPLIT distance="200" swimtime="00:03:05.87" />
                    <SPLIT distance="250" swimtime="00:03:57.87" />
                    <SPLIT distance="300" swimtime="00:04:49.92" />
                    <SPLIT distance="350" swimtime="00:05:42.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="24851" points="341" reactiontime="+108" swimtime="00:03:09.08" resultid="28245">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.45" />
                    <SPLIT distance="100" swimtime="00:01:33.54" />
                    <SPLIT distance="150" swimtime="00:02:23.47" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Carlijn" lastname="Janssen" birthdate="2010-10-14" gender="F" nation="NED" license="9256868" athleteid="28260">
              <RESULTS>
                <RESULT eventid="1053" points="610" reactiontime="+100" swimtime="00:00:26.76" resultid="28261" entrytime="00:00:28.18" entrycourse="LCM" />
                <RESULT eventid="7254" points="731" reactiontime="+94" swimtime="00:02:30.01" resultid="28262" entrytime="00:02:40.41" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.14" />
                    <SPLIT distance="100" swimtime="00:01:09.25" />
                    <SPLIT distance="150" swimtime="00:01:50.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1120" points="841" reactiontime="+85" swimtime="00:00:28.92" resultid="28263" entrytime="00:00:30.11" entrycourse="LCM" />
                <RESULT eventid="1168" points="680" reactiontime="+90" swimtime="00:01:07.25" resultid="28264" entrytime="00:01:09.35" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="7287" points="529" reactiontime="+89" swimtime="00:01:02.10" resultid="28265" entrytime="00:01:07.36" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="24851" points="603" reactiontime="+91" swimtime="00:02:28.30" resultid="28266" entrytime="00:02:39.48" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.74" />
                    <SPLIT distance="100" swimtime="00:01:08.04" />
                    <SPLIT distance="150" swimtime="00:01:49.64" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Wouter" lastname="Diepen" birthdate="2001-09-07" gender="M" nameprefix="van" nation="NED" license="9013676" athleteid="28231">
              <RESULTS>
                <RESULT eventid="1079" points="602" reactiontime="+93" swimtime="00:00:20.07" resultid="28232" entrytime="00:00:20.55" entrycourse="LCM" />
                <RESULT eventid="1127" points="660" reactiontime="+85" swimtime="00:00:23.19" resultid="28234" entrytime="00:00:23.06" entrycourse="LCM" />
                <RESULT eventid="7264" points="767" reactiontime="+99" swimtime="00:03:34.59" resultid="28235" entrytime="00:03:33.59">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:23.48" />
                    <SPLIT distance="100" swimtime="00:00:50.35" />
                    <SPLIT distance="150" swimtime="00:01:17.80" />
                    <SPLIT distance="200" swimtime="00:01:45.43" />
                    <SPLIT distance="250" swimtime="00:02:13.43" />
                    <SPLIT distance="300" swimtime="00:02:41.00" />
                    <SPLIT distance="350" swimtime="00:03:08.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1153" points="614" reactiontime="+96" swimtime="00:00:18.60" resultid="28236" entrytime="00:00:18.37" entrycourse="LCM" />
                <RESULT eventid="1175" points="808" reactiontime="+81" swimtime="00:00:49.55" resultid="28237" entrytime="00:00:49.52">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:23.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1203" points="927" reactiontime="+86" swimtime="00:03:54.72" resultid="28238" entrytime="00:03:48.89">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.38" />
                    <SPLIT distance="100" swimtime="00:00:55.48" />
                    <SPLIT distance="150" swimtime="00:01:25.06" />
                    <SPLIT distance="200" swimtime="00:01:54.91" />
                    <SPLIT distance="250" swimtime="00:02:24.75" />
                    <SPLIT distance="300" swimtime="00:02:55.21" />
                    <SPLIT distance="350" swimtime="00:03:25.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="18215" points="733" reactiontime="+100" swimtime="00:14:50.95" resultid="29464" entrytime="00:14:24.53">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:24.62" />
                    <SPLIT distance="100" swimtime="00:00:52.26" />
                    <SPLIT distance="150" swimtime="00:01:20.50" />
                    <SPLIT distance="200" swimtime="00:01:49.38" />
                    <SPLIT distance="250" swimtime="00:02:18.22" />
                    <SPLIT distance="300" swimtime="00:02:47.13" />
                    <SPLIT distance="350" swimtime="00:03:15.79" />
                    <SPLIT distance="400" swimtime="00:03:44.61" />
                    <SPLIT distance="450" swimtime="00:04:13.44" />
                    <SPLIT distance="500" swimtime="00:04:42.11" />
                    <SPLIT distance="550" swimtime="00:05:11.01" />
                    <SPLIT distance="600" swimtime="00:05:40.14" />
                    <SPLIT distance="650" swimtime="00:06:08.93" />
                    <SPLIT distance="700" swimtime="00:06:37.91" />
                    <SPLIT distance="750" swimtime="00:07:06.79" />
                    <SPLIT distance="800" swimtime="00:07:35.97" />
                    <SPLIT distance="850" swimtime="00:08:04.97" />
                    <SPLIT distance="900" swimtime="00:08:34.01" />
                    <SPLIT distance="950" swimtime="00:09:03.23" />
                    <SPLIT distance="1000" swimtime="00:09:32.19" />
                    <SPLIT distance="1050" swimtime="00:10:01.29" />
                    <SPLIT distance="1100" swimtime="00:10:30.68" />
                    <SPLIT distance="1150" swimtime="00:11:00.18" />
                    <SPLIT distance="1200" swimtime="00:11:31.86" />
                    <SPLIT distance="1250" swimtime="00:12:12.85" />
                    <SPLIT distance="1300" swimtime="00:12:51.13" />
                    <SPLIT distance="1350" swimtime="00:13:22.39" />
                    <SPLIT distance="1400" swimtime="00:13:52.82" />
                    <SPLIT distance="1450" swimtime="00:14:22.89" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Femke" lastname="Krewinkel" birthdate="1987-11-18" gender="F" nation="NED" license="9023470" athleteid="28267">
              <RESULTS>
                <RESULT eventid="1093" points="813" reactiontime="+113" swimtime="00:17:44.00" resultid="28268" entrytime="00:17:45.13" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.70" />
                    <SPLIT distance="100" swimtime="00:01:04.18" />
                    <SPLIT distance="150" swimtime="00:01:39.32" />
                    <SPLIT distance="200" swimtime="00:02:14.33" />
                    <SPLIT distance="250" swimtime="00:02:49.73" />
                    <SPLIT distance="300" swimtime="00:03:25.84" />
                    <SPLIT distance="350" swimtime="00:04:01.94" />
                    <SPLIT distance="400" swimtime="00:04:37.98" />
                    <SPLIT distance="450" swimtime="00:05:14.26" />
                    <SPLIT distance="500" swimtime="00:05:50.47" />
                    <SPLIT distance="550" swimtime="00:06:26.47" />
                    <SPLIT distance="600" swimtime="00:07:02.94" />
                    <SPLIT distance="650" swimtime="00:07:39.03" />
                    <SPLIT distance="700" swimtime="00:08:14.95" />
                    <SPLIT distance="750" swimtime="00:08:50.61" />
                    <SPLIT distance="800" swimtime="00:09:25.67" />
                    <SPLIT distance="850" swimtime="00:10:00.82" />
                    <SPLIT distance="900" swimtime="00:10:36.61" />
                    <SPLIT distance="950" swimtime="00:11:12.43" />
                    <SPLIT distance="1000" swimtime="00:11:48.33" />
                    <SPLIT distance="1050" swimtime="00:12:23.74" />
                    <SPLIT distance="1100" swimtime="00:12:59.12" />
                    <SPLIT distance="1150" swimtime="00:13:35.37" />
                    <SPLIT distance="1200" swimtime="00:14:11.60" />
                    <SPLIT distance="1250" swimtime="00:14:47.76" />
                    <SPLIT distance="1300" swimtime="00:15:23.72" />
                    <SPLIT distance="1350" swimtime="00:15:59.15" />
                    <SPLIT distance="1400" swimtime="00:16:35.31" />
                    <SPLIT distance="1450" swimtime="00:17:10.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="7254" points="760" reactiontime="+96" swimtime="00:02:26.35" resultid="28269">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.79" />
                    <SPLIT distance="100" swimtime="00:01:10.99" />
                    <SPLIT distance="150" swimtime="00:01:49.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="7278" points="837" reactiontime="+110" swimtime="00:04:30.47" resultid="28270">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.10" />
                    <SPLIT distance="100" swimtime="00:01:02.63" />
                    <SPLIT distance="150" swimtime="00:01:37.05" />
                    <SPLIT distance="200" swimtime="00:02:12.08" />
                    <SPLIT distance="250" swimtime="00:02:47.09" />
                    <SPLIT distance="300" swimtime="00:03:21.98" />
                    <SPLIT distance="350" swimtime="00:03:56.73" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jade" lastname="Arts" birthdate="2004-09-12" gender="F" nation="NED" license="9020456" athleteid="28227">
              <RESULTS>
                <RESULT eventid="1053" points="665" reactiontime="+101" swimtime="00:00:22.86" resultid="28228" entrytime="00:00:21.95" entrycourse="LCM" />
                <RESULT eventid="1147" points="811" reactiontime="+101" swimtime="00:00:20.21" resultid="28229" entrytime="00:00:19.29" />
                <RESULT eventid="1182" points="746" reactiontime="+109" swimtime="00:00:48.70" resultid="28230" entrytime="00:00:44.56" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:21.73" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luc" lastname="Ambrosius" birthdate="1975-07-24" gender="M" nation="NED" license="79269" athleteid="28226" />
            <ATHLETE firstname="Noor" lastname="Lugt" birthdate="2011-10-04" gender="F" nameprefix="van der" nation="NED" license="9255592" athleteid="28277">
              <RESULTS>
                <RESULT eventid="1053" points="498" reactiontime="+105" swimtime="00:00:28.63" resultid="28278" entrytime="00:00:30.14" entrycourse="LCM" />
                <RESULT eventid="7278" points="557" reactiontime="+87" swimtime="00:05:35.23" resultid="28279" entrytime="00:05:45.67" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.06" />
                    <SPLIT distance="100" swimtime="00:01:18.21" />
                    <SPLIT distance="150" swimtime="00:02:03.91" />
                    <SPLIT distance="200" swimtime="00:02:48.52" />
                    <SPLIT distance="250" swimtime="00:03:33.31" />
                    <SPLIT distance="300" swimtime="00:04:17.88" />
                    <SPLIT distance="350" swimtime="00:05:01.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1168" points="519" reactiontime="+96" swimtime="00:01:13.57" resultid="28280" entrytime="00:01:13.24" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1196" points="730" reactiontime="+90" swimtime="00:05:27.38" resultid="28281">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.38" />
                    <SPLIT distance="100" swimtime="00:01:18.96" />
                    <SPLIT distance="150" swimtime="00:02:01.68" />
                    <SPLIT distance="200" swimtime="00:02:45.41" />
                    <SPLIT distance="250" swimtime="00:03:27.91" />
                    <SPLIT distance="300" swimtime="00:04:10.31" />
                    <SPLIT distance="350" swimtime="00:04:52.00" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Sanne" lastname="Reichgelt" birthdate="2012-06-18" gender="F" nation="NED" license="9259813" athleteid="28291">
              <RESULTS>
                <RESULT eventid="1053" points="467" reactiontime="+143" swimtime="00:00:33.08" resultid="28292" entrytime="00:00:32.67" entrycourse="LCM" />
                <RESULT eventid="7254" points="751" reactiontime="+106" swimtime="00:02:52.87" resultid="28293">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.37" />
                    <SPLIT distance="100" swimtime="00:01:24.49" />
                    <SPLIT distance="150" swimtime="00:02:12.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1120" points="690" reactiontime="+117" swimtime="00:00:33.81" resultid="28294" entrytime="00:00:33.08" entrycourse="LCM" />
                <RESULT eventid="1168" points="622" reactiontime="+97" swimtime="00:01:15.54" resultid="28295" entrytime="00:01:18.54" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="7287" points="459" reactiontime="+100" swimtime="00:01:16.41" resultid="28296" entrytime="00:01:27.14" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.32" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="34" agetotalmin="18" gender="F">
              <RESULTS>
                <RESULT eventid="1217" reactiontime="+95" swimtime="00:04:51.85" resultid="29493" late="yes">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.72" />
                    <SPLIT distance="100" swimtime="00:00:57.88" />
                    <SPLIT distance="150" swimtime="00:01:37.46" />
                    <SPLIT distance="200" swimtime="00:02:24.54" />
                    <SPLIT distance="250" swimtime="00:03:00.96" />
                    <SPLIT distance="300" swimtime="00:03:44.74" />
                    <SPLIT distance="350" swimtime="00:04:16.02" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="28282" number="1" reactiontime="+95" />
                    <RELAYPOSITION athleteid="28239" number="2" reactiontime="+78" />
                    <RELAYPOSITION athleteid="28291" number="3" reactiontime="+56" />
                    <RELAYPOSITION athleteid="28271" number="4" reactiontime="+75" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="15" agetotalmin="14" gender="F" name="PONTOS DC" number="1">
              <RESULTS>
                <RESULT eventid="1217" reactiontime="+96" swimtime="00:04:26.28" resultid="28297" entrytime="00:04:29.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.66" />
                    <SPLIT distance="100" swimtime="00:00:56.84" />
                    <SPLIT distance="150" swimtime="00:01:30.64" />
                    <SPLIT distance="200" swimtime="00:02:10.49" />
                    <SPLIT distance="250" swimtime="00:02:40.60" />
                    <SPLIT distance="300" swimtime="00:03:16.15" />
                    <SPLIT distance="350" swimtime="00:03:48.94" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="28252" number="1" reactiontime="+96" />
                    <RELAYPOSITION athleteid="28246" number="2" reactiontime="+55" />
                    <RELAYPOSITION athleteid="28260" number="3" reactiontime="+55" />
                    <RELAYPOSITION athleteid="28277" number="4" reactiontime="+38" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="13" agetotalmin="12" gender="F" name="PONTOS DD" number="1">
              <RESULTS>
                <RESULT eventid="26758" reactiontime="+103" swimtime="00:02:00.24" resultid="28298" entrytime="00:02:00.54">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.61" />
                    <SPLIT distance="100" swimtime="00:00:57.49" />
                    <SPLIT distance="150" swimtime="00:01:31.88" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="28260" number="1" reactiontime="+103" />
                    <RELAYPOSITION athleteid="28271" number="2" reactiontime="+73" />
                    <RELAYPOSITION athleteid="28291" number="3" reactiontime="+80" />
                    <RELAYPOSITION athleteid="28277" number="4" reactiontime="+54" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="13" agemin="12" agetotalmax="-1" agetotalmin="-1" gender="X" name="PONTOS DD BM" number="1">
              <RESULTS>
                <RESULT eventid="1140" reactiontime="+92" status="EXH" swimtime="00:04:49.37" resultid="28542">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.68" />
                    <SPLIT distance="100" swimtime="00:01:08.72" />
                    <SPLIT distance="150" swimtime="00:01:47.50" />
                    <SPLIT distance="200" swimtime="00:02:31.34" />
                    <SPLIT distance="250" swimtime="00:03:05.72" />
                    <SPLIT distance="300" swimtime="00:03:42.19" />
                    <SPLIT distance="350" swimtime="00:04:13.17" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="28271" number="1" reactiontime="+92" />
                    <RELAYPOSITION athleteid="28291" number="2" reactiontime="+62" />
                    <RELAYPOSITION athleteid="28277" number="3" reactiontime="+41" />
                    <RELAYPOSITION athleteid="28260" number="4" reactiontime="+10" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="34" agemin="18" agetotalmax="-1" agetotalmin="-1" gender="X" name="PONTOS GA" number="1">
              <RESULTS>
                <RESULT eventid="1140" swimtime="00:00:00.00" resultid="28718">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="28231" number="1" />
                    <RELAYPOSITION athleteid="28252" number="2" />
                    <RELAYPOSITION athleteid="28226" number="3" />
                    <RELAYPOSITION athleteid="28227" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
          <OFFICIALS>
            <OFFICIAL officialid="4397" firstname="Michel" grade="Tijdwaarnemer" lastname="Wekking" nation="NED" />
            <OFFICIAL officialid="1523" firstname="Brenda" gender="F" grade="Tijdwaarnemer" lastname="Wekking" nation="NED" />
            <OFFICIAL officialid="21139" firstname="Lucie" gender="F" grade="Medailles" lastname="Burgers" nation="NED" />
            <OFFICIAL officialid="6668" firstname="Debbie" gender="F" grade="Medailles" lastname="Spoor" nation="NED" />
            <OFFICIAL officialid="6665" firstname="Guus" gender="M" grade="Tijdwaarnemer" lastname="Basten" nation="NED" />
            <OFFICIAL officialid="24081" firstname="Yvette" gender="F" grade="Lijnrechter" lastname="Diepen" nameprefix="van" nation="NED" />
            <OFFICIAL officialid="5283" firstname="Yvette" gender="F" grade="Tijdwaarnemer" lastname="Diepen" nameprefix="van" nation="NED" />
            <OFFICIAL officialid="29471" firstname="Luc" gender="M" grade="Tijdwaarnemer" lastname="Ambrosius" nation="NED" />
            <OFFICIAL officialid="6666" firstname="Diana" gender="F" grade="tijdwaarnemer" lastname="Basten" nation="NED" />
            <OFFICIAL officialid="21146" firstname="Ghita" gender="F" grade="Tijdwaarnemer" lastname="Puts" nation="NED" />
            <OFFICIAL officialid="6661" firstname="Yvette" gender="F" grade="Kamprechter" lastname="Diepen" nameprefix="van" nation="NED" />
            <OFFICIAL officialid="23067" firstname="Diederick" gender="M" grade="Keerpuntcommisaris" lastname="Brouwer" nation="NED" />
            <OFFICIAL officialid="3074" firstname="Stephan" gender="M" grade="Ploegleider" lastname="Steeg" nation="NED" />
            <OFFICIAL officialid="2146" firstname="Esther" gender="F" grade="Kamprechter" lastname="Vijlbrief" nation="NED" />
            <OFFICIAL officialid="29472" firstname="Yvette" gender="F" grade="voorstart" lastname="Diepen" nameprefix="van" nation="NED" />
            <OFFICIAL officialid="1509" firstname="Ruben" grade="Tijdwaarnemer (gesto" lastname="Kervel" nation="NED" />
            <OFFICIAL officialid="3088" firstname="Theo" gender="M" grade="EHBO" lastname="Cornelissen" nation="NED" />
            <OFFICIAL officialid="1538" firstname="Inge" gender="F" grade="Secretariaat" lastname="Scherpenseel" nameprefix="van" nation="NED" />
            <OFFICIAL officialid="23159" firstname="Angelique" gender="F" grade="Tijdwaarnemer" lastname="Reuver" nameprefix="de" nation="NED" />
            <OFFICIAL officialid="24078" firstname="Debbie" gender="F" grade="Keerpuntcommissaris" lastname="Spoor" nation="NED" />
            <OFFICIAL officialid="21127" firstname="Luc" gender="M" grade="Voorstart" lastname="Ambrosius" nation="NED" />
            <OFFICIAL officialid="28777" firstname="Roy" gender="M" grade="Lijnrechter" lastname="Fleuren" nation="NED" />
            <OFFICIAL officialid="2140" firstname="Monique" gender="F" grade="Voorstart" lastname="Arts" nation="NED" />
            <OFFICIAL officialid="26603" firstname="Joyce" gender="F" grade="Secretariaat" lastname="Deckwitz" nation="NED" />
            <OFFICIAL officialid="6658" firstname="Luc" gender="M" grade="Kamprechter" lastname="Ambrosius" nation="NED" />
            <OFFICIAL officialid="23645" firstname="Erik" gender="M" grade="Op- en afbouw" lastname="Arts" nation="NED" />
            <OFFICIAL officialid="23290" firstname="Debbie" gender="F" grade="Secretariaat" lastname="Spoor" nation="NED" />
          </OFFICIALS>
        </CLUB>
        <CLUB type="CLUB" code="PIRANHA" nation="NED" clubid="18180" name="ZPV Piranha">
          <OFFICIALS>
            <OFFICIAL officialid="3075" firstname="Mila" gender="F" grade="Ploegleider" lastname="Bom" nation="NED" />
          </OFFICIALS>
        </CLUB>
        <CLUB type="CLUB" code="NSF" nation="NGR" clubid="22874" name="Nigeria Swimming Federation" />
        <CLUB type="CLUB" code="SCDL" nation="GER" clubid="21975" name="SC DHfK Leipzig">
          <OFFICIALS>
            <OFFICIAL officialid="26638" firstname="David" gender="M" grade="Team Captain" lastname="Münch" nation="GER" />
            <OFFICIAL officialid="29435" firstname="Felix" gender="M" grade="Team Captain" lastname="Wahlstadt" nation="GER" />
          </OFFICIALS>
        </CLUB>
        <CLUB type="CLUB" code="NLFC" nation="GBR" clubid="22510" name="Northern Lights Finswimming Club" shortname="Northern Lights Finswimming Cl" />
        <CLUB type="CLUB" code="TSCB BRUCH" nation="GER" clubid="22880" name="TSC Bathyscaphe Bruchsal" shortname="TSC Bruchsal">
          <OFFICIALS>
            <OFFICIAL officialid="24202" firstname="Elke" gender="F" grade="Team Captain" lastname="Döring" nation="GER" />
          </OFFICIALS>
        </CLUB>
        <CLUB type="CLUB" nation="NED" clubid="18188" name="Unattached" />
        <CLUB type="CLUB" code="AQUANI" nation="BEL" clubid="22760" name="Aquani-Nivelles">
          <ATHLETES>
            <ATHLETE firstname="Arthur" lastname="Brusten" birthdate="1997-12-15" gender="M" nation="BEL" athleteid="29438">
              <RESULTS>
                <RESULT eventid="1127" points="901" reactiontime="+85" swimtime="00:00:20.91" resultid="29443" late="yes" entrytime="00:00:21.98" />
                <RESULT eventid="1175" points="998" reactiontime="+85" swimtime="00:00:46.18" resultid="29444" late="yes" entrytime="00:00:50.01">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:21.60" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lena" lastname="Druez" birthdate="2005-12-21" gender="F" nation="BEL" athleteid="29439">
              <RESULTS>
                <RESULT eventid="1120" points="792" reactiontime="+87" swimtime="00:00:25.21" resultid="29445" late="yes" entrytime="00:00:25.12" />
                <RESULT eventid="7254" points="659" reactiontime="+89" swimtime="00:02:06.97" resultid="29446" late="yes" entrytime="00:02:02.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.52" />
                    <SPLIT distance="100" swimtime="00:01:00.66" />
                    <SPLIT distance="150" swimtime="00:01:34.14" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Aloïse" lastname="Glorieuz" birthdate="2007-07-10" gender="F" nation="BEL" athleteid="29440">
              <RESULTS>
                <RESULT comment="A1 - Bewogen of te vroeg weg bij de start (geen tijd noteren)" eventid="1120" reactiontime="+73" status="DSQ" swimtime="00:00:27.73" resultid="29441" late="yes" entrytime="00:00:26.23" />
                <RESULT eventid="7254" points="681" reactiontime="+93" swimtime="00:02:15.71" resultid="29442" late="yes" entrytime="00:02:09.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.45" />
                    <SPLIT distance="100" swimtime="00:01:05.21" />
                    <SPLIT distance="150" swimtime="00:01:41.64" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <OFFICIALS>
            <OFFICIAL officialid="24795" firstname="Dominique" gender="M" grade="Team Captain" lastname="André" nation="BEL" />
          </OFFICIALS>
        </CLUB>
        <CLUB type="CLUB" code="LANAP" nation="FRA" clubid="22871" name="Longwy Apnée Nage Avec Palmes" />
        <CLUB type="CLUB" code="CSG" nation="FRA" clubid="24025" name="Club Sportif de Gravenchon" shortname="CSG">
          <ATHLETES>
            <ATHLETE firstname="Manon" lastname="Douyere" birthdate="1999-01-01" gender="F" nation="FRA" license="FRA0001060" athleteid="28477">
              <RESULTS>
                <RESULT eventid="7278" points="1141" reactiontime="+103" swimtime="00:03:34.46" resultid="28479" entrytime="00:03:30.55">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.26" />
                    <SPLIT distance="100" swimtime="00:00:53.11" />
                    <SPLIT distance="150" swimtime="00:01:20.15" />
                    <SPLIT distance="200" swimtime="00:01:47.39" />
                    <SPLIT distance="250" swimtime="00:02:14.42" />
                    <SPLIT distance="300" swimtime="00:02:41.43" />
                    <SPLIT distance="350" swimtime="00:03:08.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1147" points="1069" reactiontime="+98" swimtime="00:00:18.43" resultid="28480" entrytime="00:00:17.95" />
                <RESULT eventid="7287" points="1136" reactiontime="+103" swimtime="00:00:44.00" resultid="28481" entrytime="00:00:41.94">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:21.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="26746" points="1551" reactiontime="+132" swimtime="00:06:39.25" resultid="29434" entrytime="00:06:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:24.79" />
                    <SPLIT distance="100" swimtime="00:00:48.33" />
                    <SPLIT distance="150" swimtime="00:01:12.77" />
                    <SPLIT distance="200" swimtime="00:01:37.49" />
                    <SPLIT distance="250" swimtime="00:02:02.42" />
                    <SPLIT distance="300" swimtime="00:02:27.57" />
                    <SPLIT distance="350" swimtime="00:02:52.72" />
                    <SPLIT distance="400" swimtime="00:03:17.99" />
                    <SPLIT distance="450" swimtime="00:03:43.54" />
                    <SPLIT distance="500" swimtime="00:04:08.78" />
                    <SPLIT distance="550" swimtime="00:04:34.64" />
                    <SPLIT distance="600" swimtime="00:04:59.77" />
                    <SPLIT distance="650" swimtime="00:05:25.33" />
                    <SPLIT distance="700" swimtime="00:05:50.73" />
                    <SPLIT distance="750" swimtime="00:06:15.63" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jeanne" lastname="Daniel" birthdate="2005-01-01" gender="F" nation="FRA" license="FRA0001082" athleteid="28482">
              <RESULTS>
                <RESULT eventid="1053" points="903" reactiontime="+102" swimtime="00:00:20.65" resultid="28483" entrytime="00:00:19.75" />
                <RESULT eventid="7278" points="1095" reactiontime="+99" swimtime="00:03:37.44" resultid="28484" entrytime="00:03:36.97">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.36" />
                    <SPLIT distance="100" swimtime="00:00:53.94" />
                    <SPLIT distance="150" swimtime="00:01:22.44" />
                    <SPLIT distance="200" swimtime="00:01:50.26" />
                    <SPLIT distance="250" swimtime="00:02:17.50" />
                    <SPLIT distance="300" swimtime="00:02:44.64" />
                    <SPLIT distance="350" swimtime="00:03:11.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1147" points="1022" reactiontime="+95" swimtime="00:00:18.71" resultid="28485" entrytime="00:00:18.59" />
                <RESULT eventid="7287" points="1062" reactiontime="+97" swimtime="00:00:45.00" resultid="28486" entrytime="00:00:43.64">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:21.92" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Hugo" lastname="Meyer" birthdate="1998-01-01" gender="M" nation="FRA" license="FRA0000423" athleteid="28472">
              <RESULTS>
                <RESULT comment="B2 - Na start- en/of keerpunt meer dan 15 meter onder water gezwommen" eventid="1079" reactiontime="+84" status="DSQ" swimtime="00:00:00.00" resultid="28473" entrytime="00:00:15.78" />
                <RESULT eventid="1114" points="1352" reactiontime="+123" swimtime="00:02:54.34" resultid="28474" entrytime="00:02:52.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:20.26" />
                    <SPLIT distance="100" swimtime="00:00:41.63" />
                    <SPLIT distance="150" swimtime="00:01:03.10" />
                    <SPLIT distance="200" swimtime="00:01:24.71" />
                    <SPLIT distance="250" swimtime="00:01:46.68" />
                    <SPLIT distance="300" swimtime="00:02:09.17" />
                    <SPLIT distance="350" swimtime="00:02:32.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1153" points="1156" reactiontime="+93" swimtime="00:00:15.06" resultid="28475" entrytime="00:00:14.92" />
                <RESULT comment="A3 - De aangegeven zwemwijze niet uitgevoerd (oa duiken), A3 en B2" eventid="7295" reactiontime="+86" status="DSQ" swimtime="00:00:00.00" resultid="28476" entrytime="00:00:35.17">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:16.73" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <OFFICIALS>
            <OFFICIAL officialid="24200" firstname="Thomas" gender="M" grade="Team Captain" lastname="Chastagner" nation="FRA" />
          </OFFICIALS>
        </CLUB>
        <CLUB type="CLUB" code="STE AVERTI" nation="FRA" clubid="24717" name="SASNAP" />
        <CLUB type="CLUB" code="SCDL" nation="GER" clubid="28684" name="SC DHfK Leipzig Flossenschwimmen" shortname="SCDL">
          <ATHLETES>
            <ATHLETE firstname="Felix" lastname="Wahlstadt" birthdate="1999-07-16" gender="M" nation="GER" license="000267" athleteid="28685">
              <RESULTS>
                <RESULT eventid="1079" points="826" reactiontime="+80" swimtime="00:00:18.06" resultid="28686" entrytime="00:00:17.74" />
                <RESULT eventid="7264" points="902" reactiontime="+81" swimtime="00:03:23.33" resultid="28687" entrytime="00:03:21.86">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:22.20" />
                    <SPLIT distance="100" swimtime="00:00:47.33" />
                    <SPLIT distance="150" swimtime="00:01:12.63" />
                    <SPLIT distance="200" swimtime="00:01:38.39" />
                    <SPLIT distance="250" swimtime="00:02:04.69" />
                    <SPLIT distance="300" swimtime="00:02:31.28" />
                    <SPLIT distance="350" swimtime="00:02:57.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1153" points="727" reactiontime="+78" swimtime="00:00:17.58" resultid="28688" entrytime="00:00:16.80" />
                <RESULT eventid="24862" points="1030" reactiontime="+79" swimtime="00:01:30.99" resultid="28689" entrytime="00:01:29.72">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:20.14" />
                    <SPLIT distance="100" swimtime="00:00:43.26" />
                    <SPLIT distance="150" swimtime="00:01:06.98" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Alex Michael" lastname="Berger" birthdate="2008-08-07" gender="M" nation="GER" license="000000" athleteid="28696">
              <RESULTS>
                <RESULT eventid="7264" points="1109" reactiontime="+91" swimtime="00:03:47.48" resultid="28698" entrytime="00:03:55.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:22.75" />
                    <SPLIT distance="100" swimtime="00:00:51.33" />
                    <SPLIT distance="150" swimtime="00:01:21.37" />
                    <SPLIT distance="200" swimtime="00:01:51.64" />
                    <SPLIT distance="250" swimtime="00:02:22.34" />
                    <SPLIT distance="300" swimtime="00:02:53.15" />
                    <SPLIT distance="350" swimtime="00:03:23.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="16574" points="1244" reactiontime="+90" swimtime="00:08:03.89" resultid="28699" entrytime="00:08:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.38" />
                    <SPLIT distance="100" swimtime="00:00:56.06" />
                    <SPLIT distance="150" swimtime="00:01:28.68" />
                    <SPLIT distance="200" swimtime="00:01:58.72" />
                    <SPLIT distance="250" swimtime="00:02:30.19" />
                    <SPLIT distance="300" swimtime="00:03:02.11" />
                    <SPLIT distance="350" swimtime="00:03:34.20" />
                    <SPLIT distance="400" swimtime="00:04:06.36" />
                    <SPLIT distance="450" swimtime="00:04:36.86" />
                    <SPLIT distance="500" swimtime="00:05:07.33" />
                    <SPLIT distance="550" swimtime="00:05:38.55" />
                    <SPLIT distance="600" swimtime="00:06:09.48" />
                    <SPLIT distance="650" swimtime="00:06:39.88" />
                    <SPLIT distance="700" swimtime="00:07:10.07" />
                    <SPLIT distance="750" swimtime="00:07:38.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="7295" points="1019" reactiontime="+91" swimtime="00:00:45.14" resultid="28700" entrytime="00:00:44.82">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:21.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="24862" points="1045" reactiontime="+93" swimtime="00:01:44.18" resultid="28701" entrytime="00:01:42.60">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:22.70" />
                    <SPLIT distance="100" swimtime="00:00:50.08" />
                    <SPLIT distance="150" swimtime="00:01:18.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="18215" points="950" reactiontime="+84" swimtime="00:16:13.04" resultid="29463" entrytime="00:16:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:23.82" />
                    <SPLIT distance="100" swimtime="00:00:53.96" />
                    <SPLIT distance="150" swimtime="00:01:26.00" />
                    <SPLIT distance="200" swimtime="00:01:56.78" />
                    <SPLIT distance="250" swimtime="00:02:28.68" />
                    <SPLIT distance="300" swimtime="00:02:58.90" />
                    <SPLIT distance="350" swimtime="00:03:31.06" />
                    <SPLIT distance="400" swimtime="00:04:03.26" />
                    <SPLIT distance="450" swimtime="00:04:35.40" />
                    <SPLIT distance="500" swimtime="00:05:07.44" />
                    <SPLIT distance="550" swimtime="00:05:40.25" />
                    <SPLIT distance="600" swimtime="00:06:11.25" />
                    <SPLIT distance="650" swimtime="00:06:44.51" />
                    <SPLIT distance="700" swimtime="00:07:17.77" />
                    <SPLIT distance="750" swimtime="00:07:51.37" />
                    <SPLIT distance="800" swimtime="00:08:22.46" />
                    <SPLIT distance="850" swimtime="00:08:56.75" />
                    <SPLIT distance="900" swimtime="00:09:29.62" />
                    <SPLIT distance="950" swimtime="00:10:02.54" />
                    <SPLIT distance="1000" swimtime="00:10:36.43" />
                    <SPLIT distance="1050" swimtime="00:11:10.12" />
                    <SPLIT distance="1100" swimtime="00:11:43.46" />
                    <SPLIT distance="1150" swimtime="00:12:16.48" />
                    <SPLIT distance="1200" swimtime="00:12:51.57" />
                    <SPLIT distance="1250" swimtime="00:13:25.03" />
                    <SPLIT distance="1300" swimtime="00:14:00.49" />
                    <SPLIT distance="1350" swimtime="00:14:33.54" />
                    <SPLIT distance="1400" swimtime="00:15:03.91" />
                    <SPLIT distance="1450" swimtime="00:15:36.98" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ben Joseph" lastname="Schoodt" birthdate="2007-08-31" gender="M" nation="GER" license="002944" athleteid="28690">
              <RESULTS>
                <RESULT eventid="1079" points="1026" reactiontime="+104" swimtime="00:00:18.58" resultid="28691" entrytime="00:00:17.77" />
                <RESULT eventid="1153" points="927" reactiontime="+111" swimtime="00:00:17.38" resultid="28693" entrytime="00:00:16.81" />
                <RESULT eventid="7295" points="914" reactiontime="+93" swimtime="00:00:42.06" resultid="28694" entrytime="00:00:41.32">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:20.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="24862" points="1108" reactiontime="+99" swimtime="00:01:39.08" resultid="28695" entrytime="00:01:32.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:22.55" />
                    <SPLIT distance="100" swimtime="00:00:47.22" />
                    <SPLIT distance="150" swimtime="00:01:13.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="18215" points="827" reactiontime="+100" swimtime="00:15:05.14" resultid="29465" entrytime="00:14:38.94">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.96" />
                    <SPLIT distance="100" swimtime="00:00:54.49" />
                    <SPLIT distance="150" swimtime="00:01:24.32" />
                    <SPLIT distance="200" swimtime="00:01:54.81" />
                    <SPLIT distance="250" swimtime="00:02:25.12" />
                    <SPLIT distance="300" swimtime="00:02:54.91" />
                    <SPLIT distance="350" swimtime="00:03:25.01" />
                    <SPLIT distance="400" swimtime="00:03:55.46" />
                    <SPLIT distance="450" swimtime="00:04:25.16" />
                    <SPLIT distance="500" swimtime="00:04:55.31" />
                    <SPLIT distance="550" swimtime="00:05:25.85" />
                    <SPLIT distance="600" swimtime="00:05:55.48" />
                    <SPLIT distance="650" swimtime="00:06:25.79" />
                    <SPLIT distance="700" swimtime="00:06:55.74" />
                    <SPLIT distance="750" swimtime="00:07:25.77" />
                    <SPLIT distance="800" swimtime="00:07:55.55" />
                    <SPLIT distance="850" swimtime="00:08:25.65" />
                    <SPLIT distance="900" swimtime="00:08:56.26" />
                    <SPLIT distance="950" swimtime="00:09:26.35" />
                    <SPLIT distance="1000" swimtime="00:09:56.90" />
                    <SPLIT distance="1050" swimtime="00:10:27.71" />
                    <SPLIT distance="1100" swimtime="00:10:58.96" />
                    <SPLIT distance="1150" swimtime="00:11:29.66" />
                    <SPLIT distance="1200" swimtime="00:12:00.55" />
                    <SPLIT distance="1250" swimtime="00:12:31.54" />
                    <SPLIT distance="1300" swimtime="00:13:02.05" />
                    <SPLIT distance="1350" swimtime="00:13:32.66" />
                    <SPLIT distance="1400" swimtime="00:14:03.37" />
                    <SPLIT distance="1450" swimtime="00:14:34.64" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Kyra" lastname="Säbisch" birthdate="2008-07-25" gender="F" nation="GER" license="000000" athleteid="28713">
              <RESULTS>
                <RESULT eventid="1053" points="1073" reactiontime="+91" swimtime="00:00:20.92" resultid="28714" entrytime="00:00:21.10" />
                <RESULT eventid="7278" points="957" reactiontime="+100" swimtime="00:03:54.88" resultid="28715" entrytime="00:04:26.72">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:23.24" />
                    <SPLIT distance="100" swimtime="00:00:50.85" />
                    <SPLIT distance="150" swimtime="00:01:20.74" />
                    <SPLIT distance="200" swimtime="00:01:51.59" />
                    <SPLIT distance="250" swimtime="00:02:22.97" />
                    <SPLIT distance="300" swimtime="00:02:54.05" />
                    <SPLIT distance="350" swimtime="00:03:25.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="7287" points="1019" reactiontime="+94" swimtime="00:00:46.96" resultid="28716" entrytime="00:00:47.47">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:22.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="24851" points="940" reactiontime="+96" swimtime="00:01:48.19" resultid="28717" entrytime="00:01:49.11">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:23.99" />
                    <SPLIT distance="100" swimtime="00:00:51.46" />
                    <SPLIT distance="150" swimtime="00:01:20.28" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maiia" lastname="Horenok" birthdate="2008-05-28" gender="F" nation="GER" license="000000" athleteid="28707">
              <RESULTS>
                <RESULT eventid="1053" points="1448" reactiontime="+94" swimtime="00:00:18.93" resultid="28708" entrytime="00:00:18.97" />
                <RESULT eventid="1147" points="1219" reactiontime="+97" swimtime="00:00:17.98" resultid="28709" entrytime="00:00:17.51" />
                <RESULT eventid="7287" points="1414" reactiontime="+98" swimtime="00:00:42.10" resultid="28710" entrytime="00:00:42.46">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:20.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1182" points="1207" reactiontime="+118" swimtime="00:00:42.71" resultid="28711" entrytime="00:00:41.53">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:20.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="24851" points="1271" reactiontime="+101" swimtime="00:01:37.85" resultid="28712" entrytime="00:01:35.65">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:23.29" />
                    <SPLIT distance="100" swimtime="00:00:48.22" />
                    <SPLIT distance="150" swimtime="00:01:13.47" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Polina" lastname="Kulchytska" birthdate="2008-03-12" gender="F" nation="GER" license="000000" athleteid="28702">
              <RESULTS>
                <RESULT eventid="1093" points="867" reactiontime="+111" swimtime="00:16:10.24" resultid="28703" entrytime="00:15:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.29" />
                    <SPLIT distance="100" swimtime="00:00:59.87" />
                    <SPLIT distance="150" swimtime="00:01:32.81" />
                    <SPLIT distance="200" swimtime="00:02:06.39" />
                    <SPLIT distance="250" swimtime="00:02:40.49" />
                    <SPLIT distance="300" swimtime="00:03:13.16" />
                    <SPLIT distance="350" swimtime="00:03:46.55" />
                    <SPLIT distance="400" swimtime="00:04:19.08" />
                    <SPLIT distance="450" swimtime="00:04:52.62" />
                    <SPLIT distance="500" swimtime="00:05:26.02" />
                    <SPLIT distance="550" swimtime="00:05:58.43" />
                    <SPLIT distance="600" swimtime="00:06:30.34" />
                    <SPLIT distance="650" swimtime="00:07:03.11" />
                    <SPLIT distance="700" swimtime="00:07:35.46" />
                    <SPLIT distance="750" swimtime="00:08:07.94" />
                    <SPLIT distance="800" swimtime="00:08:40.01" />
                    <SPLIT distance="850" swimtime="00:09:13.13" />
                    <SPLIT distance="900" swimtime="00:09:46.20" />
                    <SPLIT distance="950" swimtime="00:10:18.97" />
                    <SPLIT distance="1000" swimtime="00:10:52.03" />
                    <SPLIT distance="1050" swimtime="00:11:23.70" />
                    <SPLIT distance="1100" swimtime="00:11:56.27" />
                    <SPLIT distance="1150" swimtime="00:12:28.93" />
                    <SPLIT distance="1200" swimtime="00:13:00.52" />
                    <SPLIT distance="1250" swimtime="00:13:32.98" />
                    <SPLIT distance="1300" swimtime="00:14:05.62" />
                    <SPLIT distance="1350" swimtime="00:14:38.02" />
                    <SPLIT distance="1400" swimtime="00:15:10.34" />
                    <SPLIT distance="1450" swimtime="00:15:41.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="7278" points="884" reactiontime="+117" swimtime="00:04:01.16" resultid="28704" entrytime="00:03:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.36" />
                    <SPLIT distance="100" swimtime="00:00:57.81" />
                    <SPLIT distance="150" swimtime="00:01:28.72" />
                    <SPLIT distance="200" swimtime="00:02:00.22" />
                    <SPLIT distance="250" swimtime="00:02:31.84" />
                    <SPLIT distance="300" swimtime="00:03:03.13" />
                    <SPLIT distance="350" swimtime="00:03:32.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1158" points="921" reactiontime="+129" swimtime="00:08:23.28" resultid="28705" entrytime="00:08:07.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.32" />
                    <SPLIT distance="100" swimtime="00:00:59.13" />
                    <SPLIT distance="150" swimtime="00:01:30.82" />
                    <SPLIT distance="200" swimtime="00:02:02.85" />
                    <SPLIT distance="250" swimtime="00:02:34.70" />
                    <SPLIT distance="300" swimtime="00:03:07.14" />
                    <SPLIT distance="350" swimtime="00:03:40.07" />
                    <SPLIT distance="400" swimtime="00:04:12.17" />
                    <SPLIT distance="450" swimtime="00:04:45.31" />
                    <SPLIT distance="500" swimtime="00:05:16.32" />
                    <SPLIT distance="550" swimtime="00:05:49.02" />
                    <SPLIT distance="600" swimtime="00:06:21.28" />
                    <SPLIT distance="650" swimtime="00:06:52.72" />
                    <SPLIT distance="700" swimtime="00:07:24.62" />
                    <SPLIT distance="750" swimtime="00:07:54.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1182" points="930" reactiontime="+123" swimtime="00:00:46.58" resultid="28706" entrytime="00:00:43.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:23.07" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="PAC" nation="FRA" clubid="21964" name="Palm Auray Club" />
        <CLUB type="CLUB" code="TCPR" nation="GER" clubid="22598" name="TC Preetz">
          <OFFICIALS>
            <OFFICIAL officialid="24194" firstname="Rolf" gender="M" grade="Team Captain" lastname="Blechschmidt" nation="GER" />
          </OFFICIALS>
        </CLUB>
        <CLUB type="CLUB" code="CHEM TC" nation="GER" clubid="27811" name="1. Chemnitzer Tauchverein eV" shortname="CHEMNITZER TC">
          <ATHLETES>
            <ATHLETE firstname="Marcel" lastname="Porges" birthdate="2005-01-01" gender="M" nation="GER" athleteid="27813">
              <RESULTS>
                <RESULT eventid="1079" points="907" reactiontime="+83" swimtime="00:00:17.51" resultid="28724" entrytime="00:00:17.20" />
                <RESULT eventid="1114" points="1092" reactiontime="+114" swimtime="00:03:07.20" resultid="28725" entrytime="00:03:11.34">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:20.98" />
                    <SPLIT distance="100" swimtime="00:00:43.65" />
                    <SPLIT distance="150" swimtime="00:01:07.18" />
                    <SPLIT distance="200" swimtime="00:01:31.36" />
                    <SPLIT distance="250" swimtime="00:01:55.67" />
                    <SPLIT distance="300" swimtime="00:02:19.82" />
                    <SPLIT distance="350" swimtime="00:02:44.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="16574" points="929" reactiontime="+83" swimtime="00:07:02.99" resultid="28726" entrytime="00:07:03.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:23.07" />
                    <SPLIT distance="100" swimtime="00:00:48.49" />
                    <SPLIT distance="150" swimtime="00:01:14.59" />
                    <SPLIT distance="200" swimtime="00:01:41.37" />
                    <SPLIT distance="250" swimtime="00:02:07.97" />
                    <SPLIT distance="300" swimtime="00:02:34.71" />
                    <SPLIT distance="350" swimtime="00:03:01.27" />
                    <SPLIT distance="400" swimtime="00:03:28.33" />
                    <SPLIT distance="450" swimtime="00:03:55.11" />
                    <SPLIT distance="500" swimtime="00:04:22.35" />
                    <SPLIT distance="550" swimtime="00:04:49.42" />
                    <SPLIT distance="600" swimtime="00:05:16.40" />
                    <SPLIT distance="650" swimtime="00:05:42.60" />
                    <SPLIT distance="700" swimtime="00:06:08.55" />
                    <SPLIT distance="750" swimtime="00:06:36.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1190" points="901" reactiontime="+100" swimtime="00:00:37.83" resultid="28727" entrytime="00:00:39.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:18.58" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Hans" lastname="Yannick" birthdate="2009-01-01" gender="M" nation="GER" athleteid="28720">
              <RESULTS>
                <RESULT eventid="1079" points="648" reactiontime="+93" swimtime="00:00:23.93" resultid="28728" entrytime="00:00:24.44" />
                <RESULT eventid="7264" points="840" reactiontime="+91" swimtime="00:04:09.53" resultid="28729" entrytime="00:04:14.81">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.81" />
                    <SPLIT distance="100" swimtime="00:00:55.60" />
                    <SPLIT distance="150" swimtime="00:01:28.86" />
                    <SPLIT distance="200" swimtime="00:02:01.35" />
                    <SPLIT distance="250" swimtime="00:02:34.55" />
                    <SPLIT distance="300" swimtime="00:03:08.21" />
                    <SPLIT distance="350" swimtime="00:03:41.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="16574" points="945" reactiontime="+92" swimtime="00:08:50.22" resultid="28730" entrytime="00:09:24.12">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.99" />
                    <SPLIT distance="100" swimtime="00:00:55.93" />
                    <SPLIT distance="150" swimtime="00:01:29.59" />
                    <SPLIT distance="200" swimtime="00:02:03.92" />
                    <SPLIT distance="250" swimtime="00:02:38.47" />
                    <SPLIT distance="300" swimtime="00:03:13.16" />
                    <SPLIT distance="350" swimtime="00:03:47.93" />
                    <SPLIT distance="400" swimtime="00:04:23.08" />
                    <SPLIT distance="450" swimtime="00:04:58.50" />
                    <SPLIT distance="500" swimtime="00:05:33.49" />
                    <SPLIT distance="550" swimtime="00:06:08.32" />
                    <SPLIT distance="600" swimtime="00:06:43.23" />
                    <SPLIT distance="650" swimtime="00:07:17.82" />
                    <SPLIT distance="700" swimtime="00:07:51.86" />
                    <SPLIT distance="750" swimtime="00:08:22.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="7295" points="610" reactiontime="+99" swimtime="00:00:53.55" resultid="28731" entrytime="00:00:53.67">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.09" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Angelina" lastname="Schwarzer" birthdate="2010-01-01" gender="F" nation="GER" athleteid="28722">
              <RESULTS>
                <RESULT eventid="1053" points="947" reactiontime="+93" swimtime="00:00:23.11" resultid="28736" entrytime="00:00:25.16" />
                <RESULT eventid="7278" points="1147" reactiontime="+98" swimtime="00:04:23.58" resultid="28737" entrytime="00:04:38.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.22" />
                    <SPLIT distance="100" swimtime="00:00:59.76" />
                    <SPLIT distance="150" swimtime="00:01:34.05" />
                    <SPLIT distance="200" swimtime="00:02:09.12" />
                    <SPLIT distance="250" swimtime="00:02:44.60" />
                    <SPLIT distance="300" swimtime="00:03:19.53" />
                    <SPLIT distance="350" swimtime="00:03:54.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1158" points="931" reactiontime="+104" swimtime="00:09:16.37" resultid="28738" entrytime="00:09:38.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.87" />
                    <SPLIT distance="100" swimtime="00:01:03.26" />
                    <SPLIT distance="150" swimtime="00:01:38.40" />
                    <SPLIT distance="200" swimtime="00:02:13.79" />
                    <SPLIT distance="250" swimtime="00:02:49.39" />
                    <SPLIT distance="300" swimtime="00:03:24.99" />
                    <SPLIT distance="350" swimtime="00:04:01.32" />
                    <SPLIT distance="400" swimtime="00:04:37.59" />
                    <SPLIT distance="450" swimtime="00:05:13.79" />
                    <SPLIT distance="500" swimtime="00:05:49.80" />
                    <SPLIT distance="550" swimtime="00:06:26.29" />
                    <SPLIT distance="600" swimtime="00:07:02.41" />
                    <SPLIT distance="650" swimtime="00:07:38.83" />
                    <SPLIT distance="700" swimtime="00:08:14.22" />
                    <SPLIT distance="750" swimtime="00:08:47.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="7287" points="836" reactiontime="+100" swimtime="00:00:53.30" resultid="28739" entrytime="00:00:53.16">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="24851" points="1095" reactiontime="+98" swimtime="00:02:01.59" resultid="28768" entrytime="00:02:12.98">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.84" />
                    <SPLIT distance="100" swimtime="00:00:59.30" />
                    <SPLIT distance="150" swimtime="00:01:32.29" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Hanna Maria" lastname="Nisch" birthdate="2011-01-01" gender="F" nation="GER" athleteid="28721">
              <RESULTS>
                <RESULT comment="A11 - Uitrusting voldoet niet aan de geldende eisen" eventid="1053" reactiontime="+98" status="DSQ" swimtime="00:00:00.00" resultid="28732" entrytime="00:00:26.26" />
                <RESULT eventid="7278" points="862" reactiontime="+100" swimtime="00:04:49.81" resultid="28733" entrytime="00:04:47.59">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.16" />
                    <SPLIT distance="100" swimtime="00:01:07.91" />
                    <SPLIT distance="150" swimtime="00:01:45.57" />
                    <SPLIT distance="200" swimtime="00:02:23.94" />
                    <SPLIT distance="250" swimtime="00:03:02.90" />
                    <SPLIT distance="300" swimtime="00:03:41.00" />
                    <SPLIT distance="350" swimtime="00:04:18.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1158" points="727" reactiontime="+100" swimtime="00:10:04.00" resultid="28734" entrytime="00:10:26.09">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.07" />
                    <SPLIT distance="100" swimtime="00:01:08.34" />
                    <SPLIT distance="150" swimtime="00:01:46.14" />
                    <SPLIT distance="200" swimtime="00:02:24.83" />
                    <SPLIT distance="250" swimtime="00:03:02.98" />
                    <SPLIT distance="300" swimtime="00:03:41.78" />
                    <SPLIT distance="350" swimtime="00:04:20.76" />
                    <SPLIT distance="400" swimtime="00:04:59.61" />
                    <SPLIT distance="450" swimtime="00:05:38.99" />
                    <SPLIT distance="500" swimtime="00:06:18.21" />
                    <SPLIT distance="550" swimtime="00:06:57.55" />
                    <SPLIT distance="600" swimtime="00:07:36.62" />
                    <SPLIT distance="650" swimtime="00:08:15.47" />
                    <SPLIT distance="700" swimtime="00:08:55.37" />
                    <SPLIT distance="750" swimtime="00:09:31.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="7287" points="633" reactiontime="+97" swimtime="00:00:58.50" resultid="28735" entrytime="00:01:01.11">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="24851" points="813" reactiontime="+97" swimtime="00:02:14.23" resultid="29145" entrytime="00:02:15.32">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.20" />
                    <SPLIT distance="100" swimtime="00:01:05.47" />
                    <SPLIT distance="150" swimtime="00:01:42.96" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jenny" lastname="Franke" birthdate="2008-01-01" gender="F" nation="GER" athleteid="28723">
              <RESULTS>
                <RESULT eventid="1053" points="936" reactiontime="+102" swimtime="00:00:21.89" resultid="28740" entrytime="00:00:21.92" />
                <RESULT eventid="1120" points="780" reactiontime="+89" swimtime="00:00:26.97" resultid="28741" entrytime="00:00:27.12" />
                <RESULT eventid="1147" points="712" reactiontime="+98" swimtime="00:00:21.51" resultid="28742" entrytime="00:00:19.76" />
                <RESULT eventid="7287" points="922" reactiontime="+98" swimtime="00:00:48.55" resultid="28743" entrytime="00:00:48.33">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:23.28" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <COACHES>
            <COACH firstname="Jana" gender="F" lastname="Porges" nation="GER" type="COACH" />
          </COACHES>
          <OFFICIALS>
            <OFFICIAL officialid="27812" firstname="David" gender="M" grade="Team Captain" lastname="Münch" nation="GER" />
            <OFFICIAL officialid="28803" firstname="Jana" gender="F" grade="Team Captain" lastname="Porges" nation="GER" />
          </OFFICIALS>
        </CLUB>
        <CLUB type="CLUB" code="SWISS" nation="SUI" clubid="28807" name="Swiss Team" shortname="Swiss">
          <ATHLETES>
            <ATHLETE firstname="Violante" lastname="Giuntini" birthdate="2009-01-01" gender="F" nation="SUI" license="SUSV 115062" athleteid="29063">
              <RESULTS>
                <RESULT eventid="1053" points="453" reactiontime="+106" swimtime="00:00:27.89" resultid="29069" entrytime="00:00:25.00" />
                <RESULT eventid="7254" points="812" reactiontime="+107" swimtime="00:02:15.83" resultid="29070" entrytime="00:02:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.91" />
                    <SPLIT distance="100" swimtime="00:01:04.90" />
                    <SPLIT distance="150" swimtime="00:01:41.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1147" points="391" reactiontime="+127" swimtime="00:00:26.25" resultid="29071" entrytime="00:00:24.00" />
                <RESULT eventid="1196" points="1006" reactiontime="+112" swimtime="00:04:43.67" resultid="29072" entrytime="00:04:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.17" />
                    <SPLIT distance="100" swimtime="00:01:05.37" />
                    <SPLIT distance="150" swimtime="00:01:41.86" />
                    <SPLIT distance="200" swimtime="00:02:18.37" />
                    <SPLIT distance="250" swimtime="00:02:56.04" />
                    <SPLIT distance="300" swimtime="00:03:33.76" />
                    <SPLIT distance="350" swimtime="00:04:09.35" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ariel" lastname="Scaglia" birthdate="2010-01-01" gender="F" nation="SUI" license="SUSV 115064" athleteid="29062">
              <RESULTS>
                <RESULT eventid="1120" points="1060" reactiontime="+87" swimtime="00:00:26.77" resultid="29074" entrytime="00:00:25.00" />
                <RESULT eventid="1168" points="974" reactiontime="+87" swimtime="00:00:59.66" resultid="29075" entrytime="00:01:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="7287" points="673" reactiontime="+86" swimtime="00:00:57.31" resultid="29076" entrytime="00:00:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1053" points="851" reactiontime="+98" swimtime="00:00:23.95" resultid="29081" entrytime="00:00:23.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lea" lastname="Del Ponte" birthdate="2005-01-01" gender="F" nation="SUI" license="SUSV 114143" athleteid="29064">
              <RESULTS>
                <RESULT eventid="1053" points="820" reactiontime="+86" swimtime="00:00:21.32" resultid="29065" entrytime="00:00:21.12" />
                <RESULT eventid="1120" points="866" reactiontime="+83" swimtime="00:00:24.47" resultid="29066" entrytime="00:00:26.00" />
                <RESULT eventid="1147" points="918" reactiontime="+98" swimtime="00:00:19.39" resultid="29067" entrytime="00:00:19.08" />
                <RESULT eventid="7287" points="898" reactiontime="+82" swimtime="00:00:47.58" resultid="29068" entrytime="00:00:47.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:21.75" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Filip" lastname="Jancev" birthdate="2009-01-01" gender="M" nation="SUI" license="SUSV 114764" athleteid="29061">
              <RESULTS>
                <RESULT eventid="7271" points="740" reactiontime="+85" swimtime="00:02:05.39" resultid="29077" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.73" />
                    <SPLIT distance="100" swimtime="00:00:57.52" />
                    <SPLIT distance="150" swimtime="00:01:31.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1175" points="790" reactiontime="+93" swimtime="00:00:54.54" resultid="29078" entrytime="00:00:56.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1127" points="767" reactiontime="+93" swimtime="00:00:24.98" resultid="29079" entrytime="00:00:24.00" />
                <RESULT eventid="1203" points="10871" reactiontime="+90" swimtime="00:04:30.84" resultid="29080" entrytime="00:04:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.32" />
                    <SPLIT distance="100" swimtime="00:00:59.36" />
                    <SPLIT distance="150" swimtime="00:01:34.05" />
                    <SPLIT distance="200" swimtime="00:02:10.62" />
                    <SPLIT distance="250" swimtime="00:02:46.66" />
                    <SPLIT distance="300" swimtime="00:03:22.83" />
                    <SPLIT distance="350" swimtime="00:03:59.22" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <OFFICIALS>
            <OFFICIAL officialid="29436" firstname="Desire" gender="F" grade="Team Captain" lastname="Tiu" nation="SUI" />
            <OFFICIAL officialid="28816" firstname="Dimitri" gender="M" grade="Team Captain" lastname="Kalas" nation="SUI" />
          </OFFICIALS>
        </CLUB>
        <CLUB type="CLUB" code="CCNAP" nation="FRA" clubid="24421" name="Club Ciotaden de Nage avec Palmes" shortname="Ciotaden NP">
          <ATHLETES>
            <ATHLETE firstname="Antonin" lastname="Lebeau" birthdate="2007-01-01" gender="M" nation="FRA" license="A-19-841353" athleteid="28851">
              <RESULTS>
                <RESULT eventid="1079" points="925" reactiontime="+93" swimtime="00:00:19.23" resultid="28852" entrytime="00:00:19.00" />
                <RESULT eventid="7264" points="1228" reactiontime="+95" swimtime="00:03:16.08" resultid="28853" entrytime="00:03:19.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:22.37" />
                    <SPLIT distance="100" swimtime="00:00:46.83" />
                    <SPLIT distance="150" swimtime="00:01:11.74" />
                    <SPLIT distance="200" swimtime="00:01:36.62" />
                    <SPLIT distance="250" swimtime="00:02:01.70" />
                    <SPLIT distance="300" swimtime="00:02:26.89" />
                    <SPLIT distance="350" swimtime="00:02:51.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="16574" points="1278" reactiontime="+97" swimtime="00:06:50.52" resultid="28854" entrytime="00:06:53.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:21.92" />
                    <SPLIT distance="100" swimtime="00:00:46.00" />
                    <SPLIT distance="150" swimtime="00:01:10.90" />
                    <SPLIT distance="200" swimtime="00:01:36.27" />
                    <SPLIT distance="250" swimtime="00:02:02.19" />
                    <SPLIT distance="300" swimtime="00:02:28.21" />
                    <SPLIT distance="350" swimtime="00:02:54.15" />
                    <SPLIT distance="400" swimtime="00:03:20.48" />
                    <SPLIT distance="450" swimtime="00:03:46.61" />
                    <SPLIT distance="500" swimtime="00:04:12.73" />
                    <SPLIT distance="550" swimtime="00:04:39.15" />
                    <SPLIT distance="600" swimtime="00:05:05.72" />
                    <SPLIT distance="650" swimtime="00:05:31.90" />
                    <SPLIT distance="700" swimtime="00:05:58.51" />
                    <SPLIT distance="750" swimtime="00:06:24.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="24862" points="1399" reactiontime="+97" swimtime="00:01:31.68" resultid="28855" entrytime="00:01:30.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:21.30" />
                    <SPLIT distance="100" swimtime="00:00:44.43" />
                    <SPLIT distance="150" swimtime="00:01:07.87" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <OFFICIALS>
            <OFFICIAL officialid="24482" firstname="Benoit" gender="M" grade="Team Captain" lastname="Lebeau" nation="FRA" />
            <OFFICIAL officialid="24420" firstname="Jean Marc" gender="M" grade="Team Captain" lastname="Perkovic" nation="FRA" />
          </OFFICIALS>
        </CLUB>
        <CLUB type="CLUB" code="WAVES" nation="NED" clubid="26791" name="Waves" shortname="Vinzwemvereniging WAVES">
          <ATHLETES>
            <ATHLETE firstname="Mette" lastname="Munk" birthdate="2005-04-24" gender="F" nameprefix="de" nation="NED" license="9024160" athleteid="28184" level="A/B/C">
              <RESULTS>
                <RESULT eventid="1053" points="534" reactiontime="+121" swimtime="00:00:24.60" resultid="28185" />
                <RESULT eventid="7254" points="628" reactiontime="+92" swimtime="00:02:09.07" resultid="28186" entrytime="00:02:17.46" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.45" />
                    <SPLIT distance="100" swimtime="00:01:01.76" />
                    <SPLIT distance="150" swimtime="00:01:35.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1120" points="611" reactiontime="+96" swimtime="00:00:27.48" resultid="28187" />
                <RESULT eventid="1168" points="618" reactiontime="+93" swimtime="00:00:59.63" resultid="28188" entrytime="00:01:01.61" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1196" points="787" reactiontime="+101" swimtime="00:04:45.94" resultid="28189" entrytime="00:05:05.72" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.02" />
                    <SPLIT distance="100" swimtime="00:01:07.13" />
                    <SPLIT distance="150" swimtime="00:01:43.96" />
                    <SPLIT distance="200" swimtime="00:02:20.98" />
                    <SPLIT distance="250" swimtime="00:02:58.77" />
                    <SPLIT distance="300" swimtime="00:03:36.20" />
                    <SPLIT distance="350" swimtime="00:04:13.48" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Richard" lastname="Peters" birthdate="2004-06-23" gender="M" nation="NED" license="9028312" athleteid="28190">
              <RESULTS>
                <RESULT comment="B2 - Na start- en/of keerpunt meer dan 15 meter onder water gezwommen" eventid="1079" reactiontime="+96" status="DSQ" swimtime="00:00:22.13" resultid="28191" />
                <RESULT eventid="7271" points="778" reactiontime="+91" swimtime="00:01:58.48" resultid="28192">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.02" />
                    <SPLIT distance="100" swimtime="00:00:56.92" />
                    <SPLIT distance="150" swimtime="00:01:27.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1127" points="541" reactiontime="+95" swimtime="00:00:24.78" resultid="28193" />
                <RESULT eventid="1153" points="448" reactiontime="+92" swimtime="00:00:20.66" resultid="28194" />
                <RESULT eventid="7295" points="493" reactiontime="+101" swimtime="00:00:49.88" resultid="28195">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:23.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="24862" points="522" reactiontime="+95" swimtime="00:01:54.13" resultid="28196">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:24.35" />
                    <SPLIT distance="100" swimtime="00:00:52.60" />
                    <SPLIT distance="150" swimtime="00:01:23.79" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marco" lastname="Rutten" birthdate="1971-09-05" gender="M" nation="NED" license="9261638" athleteid="28204">
              <RESULTS>
                <RESULT eventid="1079" points="751" reactiontime="+101" swimtime="00:00:23.38" resultid="28205" entrytime="00:00:23.83" entrycourse="LCM" />
                <RESULT eventid="7271" points="815" reactiontime="+98" swimtime="00:02:05.86" resultid="28206" entrytime="00:02:06.25" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.85" />
                    <SPLIT distance="100" swimtime="00:00:58.73" />
                    <SPLIT distance="150" swimtime="00:01:32.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1127" points="737" reactiontime="+99" swimtime="00:00:25.34" resultid="28207" entrytime="00:00:25.10" entrycourse="LCM" />
                <RESULT eventid="1153" points="644" reactiontime="+103" swimtime="00:00:21.44" resultid="28208" entrytime="00:00:21.93" entrycourse="LCM" />
                <RESULT eventid="1175" points="807" reactiontime="+94" swimtime="00:00:55.74" resultid="28209" entrytime="00:00:56.44" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.69" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Nederlands record" eventid="1203" points="1000" reactiontime="+95" swimtime="00:04:44.84" resultid="28210">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.52" />
                    <SPLIT distance="100" swimtime="00:01:03.48" />
                    <SPLIT distance="150" swimtime="00:01:37.95" />
                    <SPLIT distance="200" swimtime="00:02:14.06" />
                    <SPLIT distance="250" swimtime="00:02:50.46" />
                    <SPLIT distance="300" swimtime="00:03:28.57" />
                    <SPLIT distance="350" swimtime="00:04:07.89" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Isa" lastname="Rutten" birthdate="2004-05-12" gender="F" nation="NED" license="9218514" athleteid="28197">
              <RESULTS>
                <RESULT eventid="1053" points="479" reactiontime="+113" swimtime="00:00:25.50" resultid="28198" entrytime="00:00:24.87" entrycourse="LCM" />
                <RESULT eventid="7254" points="547" reactiontime="+94" swimtime="00:02:15.13" resultid="28199" entrytime="00:02:16.42" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.36" />
                    <SPLIT distance="100" swimtime="00:01:05.66" />
                    <SPLIT distance="150" swimtime="00:01:41.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1120" points="585" reactiontime="+96" swimtime="00:00:27.89" resultid="28200" entrytime="00:00:26.74" entrycourse="LCM" />
                <RESULT eventid="1147" points="387" reactiontime="+110" swimtime="00:00:25.85" resultid="28201" entrytime="00:00:24.71" entrycourse="LCM" />
                <RESULT eventid="1168" points="593" reactiontime="+92" swimtime="00:01:00.46" resultid="28202" entrytime="00:01:01.84" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="7287" points="521" reactiontime="+107" swimtime="00:00:57.04" resultid="28203" entrytime="00:00:56.76" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.89" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Allard" lastname="Wagensveld" birthdate="1974-05-30" gender="M" nation="NED" license="9024164" athleteid="28218">
              <RESULTS>
                <RESULT eventid="1079" points="671" reactiontime="+102" swimtime="00:00:21.78" resultid="28219" entrytime="00:00:21.84" entrycourse="LCM" />
                <RESULT eventid="7271" points="807" reactiontime="+94" swimtime="00:02:03.72" resultid="28220" entrytime="00:02:03.78" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.84" />
                    <SPLIT distance="100" swimtime="00:00:57.07" />
                    <SPLIT distance="150" swimtime="00:01:29.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1127" points="810" reactiontime="+90" swimtime="00:00:24.26" resultid="28221" entrytime="00:00:24.26" entrycourse="LCM" />
                <RESULT eventid="1153" points="813" reactiontime="+112" swimtime="00:00:19.41" resultid="28222" entrytime="00:00:19.49" entrycourse="LCM" />
                <RESULT eventid="1175" points="843" reactiontime="+96" swimtime="00:00:53.56" resultid="28223" entrytime="00:00:53.56" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="7295" points="854" reactiontime="+97" swimtime="00:00:47.86" resultid="28224" entrytime="00:00:48.38" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:23.41" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Nederlands record" eventid="1190" points="1135" reactiontime="+126" swimtime="00:00:45.50" resultid="28225" entrytime="00:00:47.26" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:22.21" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Sije" lastname="Veenstra" birthdate="2006-09-24" gender="M" nation="NED" license="9258112" athleteid="28211">
              <RESULTS>
                <RESULT eventid="1079" points="365" reactiontime="+109" swimtime="00:00:26.21" resultid="28212" />
                <RESULT eventid="7271" points="572" reactiontime="+106" swimtime="00:02:15.41" resultid="28213">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.23" />
                    <SPLIT distance="100" swimtime="00:01:02.26" />
                    <SPLIT distance="150" swimtime="00:01:38.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1127" points="587" reactiontime="+109" swimtime="00:00:27.00" resultid="28214" />
                <RESULT eventid="1175" points="622" reactiontime="+103" swimtime="00:00:58.80" resultid="28215">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="7295" points="351" reactiontime="+99" swimtime="00:00:57.84" resultid="28216">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="24862" points="421" reactiontime="+110" swimtime="00:02:16.75" resultid="28217">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.60" />
                    <SPLIT distance="100" swimtime="00:01:03.84" />
                    <SPLIT distance="150" swimtime="00:01:40.43" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Coen" lastname="Bronkhorst" birthdate="2004-04-08" gender="M" nation="NED" license="9021604" athleteid="28178">
              <RESULTS>
                <RESULT eventid="1079" points="489" reactiontime="+119" swimtime="00:00:21.50" resultid="28179" entrytime="00:00:21.87" entrycourse="LCM" />
                <RESULT eventid="7271" points="751" reactiontime="+95" swimtime="00:01:59.87" resultid="28180" entrytime="00:01:59.86" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.06" />
                    <SPLIT distance="100" swimtime="00:00:58.86" />
                    <SPLIT distance="150" swimtime="00:01:30.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1127" points="576" reactiontime="+98" swimtime="00:00:24.27" resultid="28181" entrytime="00:00:23.76" entrycourse="LCM" />
                <RESULT eventid="7295" points="564" reactiontime="+118" swimtime="00:00:47.70" resultid="28182" entrytime="00:00:50.43" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:23.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="24862" points="367" reactiontime="+120" swimtime="00:02:08.34" resultid="28183" entrytime="00:02:04.99" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.80" />
                    <SPLIT distance="100" swimtime="00:01:00.81" />
                    <SPLIT distance="150" swimtime="00:01:34.89" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="34" agetotalmin="18" gender="M" name="WAVES HA" number="1">
              <RESULTS>
                <RESULT eventid="26768" reactiontime="+103" swimtime="00:01:35.88" resultid="29481">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:24.85" />
                    <SPLIT distance="100" swimtime="00:00:52.16" />
                    <SPLIT distance="150" swimtime="00:01:14.26" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="28204" number="1" reactiontime="+103" />
                    <RELAYPOSITION athleteid="28211" number="2" reactiontime="+61" />
                    <RELAYPOSITION athleteid="28218" number="3" reactiontime="+38" />
                    <RELAYPOSITION athleteid="28178" number="4" reactiontime="+40" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="34" agetotalmin="18" gender="M" name="WAVES HA" number="1">
              <RESULTS>
                <RESULT eventid="24873" reactiontime="+99" swimtime="00:03:18.97" resultid="29484">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.58" />
                    <SPLIT distance="100" swimtime="00:00:53.47" />
                    <SPLIT distance="150" swimtime="00:01:16.91" />
                    <SPLIT distance="200" swimtime="00:01:42.75" />
                    <SPLIT distance="250" swimtime="00:02:06.63" />
                    <SPLIT distance="300" swimtime="00:02:30.93" />
                    <SPLIT distance="350" swimtime="00:02:53.93" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="28204" number="1" reactiontime="+99" />
                    <RELAYPOSITION athleteid="28190" number="2" reactiontime="+29" />
                    <RELAYPOSITION athleteid="28178" number="3" reactiontime="+68" />
                    <RELAYPOSITION athleteid="28218" number="4" reactiontime="+44" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="34" agemin="18" agetotalmax="-1" agetotalmin="-1" gender="X" name="Waves GA" number="1">
              <RESULTS>
                <RESULT comment="Nederlands record" eventid="1140" reactiontime="+93" swimtime="00:03:49.47" resultid="29482">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.80" />
                    <SPLIT distance="100" swimtime="00:00:54.06" />
                    <SPLIT distance="150" swimtime="00:01:24.76" />
                    <SPLIT distance="200" swimtime="00:01:56.74" />
                    <SPLIT distance="250" swimtime="00:02:25.07" />
                    <SPLIT distance="300" swimtime="00:02:57.09" />
                    <SPLIT distance="350" swimtime="00:03:22.36" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="28178" number="1" reactiontime="+93" />
                    <RELAYPOSITION athleteid="28197" number="2" reactiontime="+44" />
                    <RELAYPOSITION athleteid="28184" number="3" reactiontime="+13" />
                    <RELAYPOSITION athleteid="28190" number="4" reactiontime="+36" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="34" agetotalmin="18" gender="X" name="WAVES GA" number="1">
              <RESULTS>
                <RESULT eventid="1210" reactiontime="+98" swimtime="00:01:28.72" resultid="29483">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:20.30" />
                    <SPLIT distance="100" swimtime="00:00:43.67" />
                    <SPLIT distance="150" swimtime="00:01:09.00" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="28190" number="1" reactiontime="+98" />
                    <RELAYPOSITION athleteid="28184" number="2" />
                    <RELAYPOSITION athleteid="28197" number="3" />
                    <RELAYPOSITION athleteid="28178" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
          <OFFICIALS>
            <OFFICIAL officialid="25528" firstname="Joyce" gender="F" grade="Tijdwaarnemer" lastname="Giessen" nameprefix="van der" nation="NED" />
            <OFFICIAL officialid="27676" firstname="Els" gender="F" grade="Ploegleider" lastname="Smilde" nation="NED" />
            <OFFICIAL officialid="18262" firstname="Mirjam" gender="F" grade="Tijdwaarnemer" lastname="Munk" nameprefix="de" nation="NED" />
          </OFFICIALS>
        </CLUB>
        <CLUB type="CLUB" code="SSC HALLE" nation="GER" clubid="27900" name="SSC Halle">
          <OFFICIALS>
            <OFFICIAL officialid="27902" firstname="Jörg" gender="M" grade="Team Captain" lastname="Hoffman" nation="GER" />
          </OFFICIALS>
        </CLUB>
        <CLUB type="UNATTACHED">
          <OFFICIALS>
            <OFFICIAL officialid="21136" firstname="John" gender="M" grade="Medailles" lastname="Schokx" />
            <OFFICIAL officialid="3086" firstname="Hylke" grade="Speaker" lastname="Faas" />
            <OFFICIAL officialid="18251" firstname="Evert" gender="M" grade="Tijdwaarnemer" lastname="Calor" />
            <OFFICIAL officialid="26602" firstname="Arien" gender="M" grade="Elec. Tijdwaarneming" lastname="Korte" nameprefix="de" />
            <OFFICIAL officialid="18264" firstname="Günter" gender="M" grade="Tijdwaarnemer" lastname="Käseberg" />
            <OFFICIAL officialid="26601" firstname="Kees Jan" gender="M" grade="Elec. Tijdwaarneming" lastname="Dijk" nameprefix="van" />
            <OFFICIAL officialid="21145" firstname="Hélène" gender="F" grade="Coörd. Estafettes" lastname="Bouwmeester" />
            <OFFICIAL officialid="24077" firstname="Hans" gender="M" grade="Keerpuntcommissaris" lastname="Liefland" nameprefix="van" />
            <OFFICIAL officialid="7483" firstname="Bijspringen recordaanvragen" grade="tijdwaarnemer" lastname="Diederick, Marc, Dick" />
            <OFFICIAL officialid="18261" />
            <OFFICIAL officialid="21141" firstname="Joris" gender="M" grade="Video opnames" lastname="Robijn" />
            <OFFICIAL officialid="2150" gender="F" grade="Speaker" lastname="SPEAKER" />
            <OFFICIAL officialid="25529" firstname="Heike" gender="F" grade="Tijdwaarnemer" lastname="Bieler" />
            <OFFICIAL officialid="26637" gender="M" />
            <OFFICIAL officialid="28783" firstname="Manfred" gender="M" grade="Tijdwaarnemer" lastname="Jöckel" />
            <OFFICIAL officialid="21317" firstname="Marleen" gender="F" grade="Voorstart" lastname="Enter" />
            <OFFICIAL officialid="18242" firstname="Jan" gender="M" grade="Elec. Tijdwaarneming" lastname="Ven" nameprefix="van de" />
            <OFFICIAL officialid="24187" firstname="Via Karin" gender="M" lastname="OVERIGE INDELING " />
            <OFFICIAL officialid="18254" firstname="Free" gender="M" grade="Lijnrechter" lastname="Deurinxk" />
          </OFFICIALS>
        </CLUB>
      </CLUBS>
    </MEET>
  </MEETS>
  <TIMESTANDARDLISTS>
    <TIMESTANDARDLIST timestandardlistid="3540" course="LCM" gender="M" name="Vinzwemmen tijdstandaarden" type="DEFAULT">
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:00:03.30">
          <SWIMSTYLE distance="25" relaycount="1" stroke="BIFINS" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:19.00">
          <SWIMSTYLE distance="1500" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:02.30">
          <SWIMSTYLE distance="100" relaycount="1" stroke="IMMERSION" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:05.30">
          <SWIMSTYLE distance="400" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:07.00">
          <SWIMSTYLE distance="100" relaycount="4" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:03.30">
          <SWIMSTYLE distance="200" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:02.00">
          <SWIMSTYLE distance="25" relaycount="1" stroke="BIFINS" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:05.30">
          <SWIMSTYLE distance="400" relaycount="1" stroke="IMMERSION" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:10.00">
          <SWIMSTYLE distance="800" relaycount="1" stroke="IMMERSION" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:02.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="APNEA" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:11.00">
          <SWIMSTYLE distance="800" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:12.00">
          <SWIMSTYLE distance="200" relaycount="4" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:02.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:02.30">
          <SWIMSTYLE distance="100" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:02.00">
          <SWIMSTYLE distance="25" relaycount="1" stroke="BIFINS" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="3541" course="SCM" gender="M" name="Vinzwemmen tijdstandaarden" type="DEFAULT">
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:00:19.00">
          <SWIMSTYLE distance="1500" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:02.30">
          <SWIMSTYLE distance="100" relaycount="1" stroke="IMMERSION" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:05.30">
          <SWIMSTYLE distance="400" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:07.00">
          <SWIMSTYLE distance="100" relaycount="4" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:03.30">
          <SWIMSTYLE distance="200" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:05.30">
          <SWIMSTYLE distance="400" relaycount="1" stroke="IMMERSION" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:02.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="APNEA" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:11.00">
          <SWIMSTYLE distance="800" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:12.00">
          <SWIMSTYLE distance="200" relaycount="4" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:02.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:02.30">
          <SWIMSTYLE distance="100" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="3542" course="LCM" gender="F" name="Vinzwemmen tijdstandaarden" type="DEFAULT">
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:00:03.30">
          <SWIMSTYLE distance="25" relaycount="1" stroke="BIFINS" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:19.00">
          <SWIMSTYLE distance="1500" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:02.30">
          <SWIMSTYLE distance="100" relaycount="1" stroke="IMMERSION" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:05.30">
          <SWIMSTYLE distance="400" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:07.00">
          <SWIMSTYLE distance="100" relaycount="4" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:03.30">
          <SWIMSTYLE distance="200" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:02.00">
          <SWIMSTYLE distance="25" relaycount="1" stroke="BIFINS" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:05.30">
          <SWIMSTYLE distance="400" relaycount="1" stroke="IMMERSION" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:10.00">
          <SWIMSTYLE distance="800" relaycount="1" stroke="IMMERSION" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:02.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="APNEA" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:11.00">
          <SWIMSTYLE distance="800" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:12.00">
          <SWIMSTYLE distance="200" relaycount="4" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:02.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:02.30">
          <SWIMSTYLE distance="100" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:02.00">
          <SWIMSTYLE distance="25" relaycount="1" stroke="BIFINS" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="3543" course="SCM" gender="F" name="Vinzwemmen tijdstandaarden" type="DEFAULT">
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:00:19.00">
          <SWIMSTYLE distance="1500" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:02.30">
          <SWIMSTYLE distance="100" relaycount="1" stroke="IMMERSION" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:05.30">
          <SWIMSTYLE distance="400" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:07.00">
          <SWIMSTYLE distance="100" relaycount="4" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:03.30">
          <SWIMSTYLE distance="200" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:05.30">
          <SWIMSTYLE distance="400" relaycount="1" stroke="IMMERSION" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:02.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="APNEA" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:11.00">
          <SWIMSTYLE distance="800" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:12.00">
          <SWIMSTYLE distance="200" relaycount="4" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:02.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:02.30">
          <SWIMSTYLE distance="100" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
  </TIMESTANDARDLISTS>
</LENEX>
