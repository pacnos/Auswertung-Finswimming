<?xml version="1.0" encoding="UTF-8"?>
<LENEX version="3.0">
  <CONSTRUCTOR name="EasyWk" version="5.23 BETA" registration="">
    <CONTACT name="Bjoern Stickan" internet="http://www.easywk.de" email="info@easywk.de" />
  </CONSTRUCTOR>
  <MEETS>
    <MEET city="Zwickau" course="LCM" name="33. offene Sachsenmeisterschaften und 16. Sachsenmeisterschaften der Masters im Finswimming" nation="GER" organizer="TC Manta Zwickau e.V." hostclub="Landestauchsportverband Sachsen e.V." deadline="2023-03-23" timing="AUTOMATIC">
      <CONTACT city="Leipzig" email="sachsenmeisterschaften@egd-tb.de" fax="+49 (0) 341 4426911" name="Brandenburg, Thilo" phone="+49 (0) 178 8150839" street="Zum Leutzscher Holz 26" zip="04178" />
      <AGEDATE type="YEAR" value="2023-01-01" />
      <SESSIONS>
        <SESSION number="1" date="2023-04-01" daytime="09:20" officialmeeting="08:30" warmupfrom="08:00">
          <EVENTS>
            <EVENT eventid="1" number="1" gender="F" round="TIM">
              <SWIMSTYLE stroke="SURFACE" relaycount="1" distance="400" />
              <FEE value="600" currency="EUR" />
              <HEATS>
                <HEAT heatid="1001" number="1" />
                <HEAT heatid="1002" number="2" />
                <HEAT heatid="1003" number="3" />
                <HEAT heatid="1004" number="4" />
                <HEAT heatid="1005" number="5" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="10" agemin="7" name="Sachsen - Altersklasse F" />
                <AGEGROUP agegroupid="2" agemax="11" agemin="11" name="Sachsen - Altersklasse E">
                  <RANKINGS>
                    <RANKING place="1" resultid="347" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3" agemax="13" agemin="12" name="Sachsen - Altersklasse D">
                  <RANKINGS>
                    <RANKING place="1" resultid="280" />
                    <RANKING place="4" resultid="291" />
                    <RANKING place="5" resultid="375" />
                    <RANKING place="6" resultid="393" />
                    <RANKING place="3" resultid="397" />
                    <RANKING place="2" resultid="490" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="15" agemin="14" name="Sachsen - Altersklasse C">
                  <RANKINGS>
                    <RANKING place="1" resultid="470" />
                    <RANKING place="2" resultid="706" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="17" agemin="16" name="Sachsen - Altersklasse B">
                  <RANKINGS>
                    <RANKING place="1" resultid="464" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6" agemax="34" agemin="18" name="Sachsen - Altersklasse A">
                  <RANKINGS>
                    <RANKING place="4" resultid="413" />
                    <RANKING place="1" resultid="487" />
                    <RANKING place="3" resultid="635" />
                    <RANKING place="2" resultid="652" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7" agemax="10" agemin="7" name="offen - Altersklasse F">
                  <RANKINGS>
                    <RANKING place="1" resultid="100" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8" agemax="11" agemin="11" name="offen - Altersklasse E">
                  <RANKINGS>
                    <RANKING place="1" resultid="347" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9" agemax="13" agemin="12" name="offen - Altersklasse D">
                  <RANKINGS>
                    <RANKING place="7" resultid="93" />
                    <RANKING place="1" resultid="280" />
                    <RANKING place="4" resultid="291" />
                    <RANKING place="5" resultid="375" />
                    <RANKING place="6" resultid="393" />
                    <RANKING place="3" resultid="397" />
                    <RANKING place="2" resultid="490" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10" agemax="15" agemin="14" name="offen - Altersklasse C">
                  <RANKINGS>
                    <RANKING place="1" resultid="470" />
                    <RANKING place="2" resultid="556" />
                    <RANKING place="4" resultid="693" />
                    <RANKING place="3" resultid="706" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11" agemax="17" agemin="16" name="offen - Altersklasse B">
                  <RANKINGS>
                    <RANKING place="3" resultid="12" />
                    <RANKING place="1" resultid="65" />
                    <RANKING place="4" resultid="251" />
                    <RANKING place="5" resultid="464" />
                    <RANKING place="2" resultid="561" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="12" agemax="34" agemin="18" name="offen - Altersklasse A">
                  <RANKINGS>
                    <RANKING place="6" resultid="27" />
                    <RANKING place="5" resultid="110" />
                    <RANKING place="7" resultid="413" />
                    <RANKING place="2" resultid="487" />
                    <RANKING place="1" resultid="543" />
                    <RANKING place="4" resultid="635" />
                    <RANKING place="3" resultid="652" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="13" agemax="44" agemin="35" name="Sachsen - Masters AK I">
                  <RANKINGS>
                    <RANKING place="1" resultid="604" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="14" agemax="45" agemin="36" name="Sachsen - Masters AK II">
                  <RANKINGS>
                    <RANKING place="1" resultid="604" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15" agemax="55" agemin="46" name="Sachsen - Masters AK III" />
                <AGEGROUP agegroupid="16" agemax="65" agemin="56" name="Sachsen - Masters AK IV" />
                <AGEGROUP agegroupid="17" agemax="-1" agemin="66" name="Sachsen - Masters AK V" />
                <AGEGROUP agegroupid="18" agemax="44" agemin="35" name="offen - Masters AK I">
                  <RANKINGS>
                    <RANKING place="1" resultid="604" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="19" agemax="45" agemin="36" name="offen - Masters AK II">
                  <RANKINGS>
                    <RANKING place="1" resultid="604" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="20" agemax="55" agemin="46" name="offen - Masters AK III">
                  <RANKINGS>
                    <RANKING place="1" resultid="197" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="21" agemax="65" agemin="56" name="offen - Masters AK IV">
                  <RANKINGS>
                    <RANKING place="1" resultid="699" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="22" agemax="-1" agemin="66" name="offen - Masters AK V" />
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="2" number="2" gender="M" round="TIM">
              <SWIMSTYLE stroke="SURFACE" relaycount="1" distance="400" />
              <FEE value="600" currency="EUR" />
              <HEATS>
                <HEAT heatid="2001" number="1" />
                <HEAT heatid="2002" number="2" />
                <HEAT heatid="2003" number="3" />
                <HEAT heatid="2004" number="4" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="10" agemin="7" name="Sachsen - Altersklasse F">
                  <RANKINGS>
                    <RANKING place="1" resultid="273" />
                    <RANKING place="2" resultid="329" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2" agemax="11" agemin="11" name="Sachsen - Altersklasse E" />
                <AGEGROUP agegroupid="3" agemax="13" agemin="12" name="Sachsen - Altersklasse D" />
                <AGEGROUP agegroupid="4" agemax="15" agemin="14" name="Sachsen - Altersklasse C">
                  <RANKINGS>
                    <RANKING place="1" resultid="433" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="17" agemin="16" name="Sachsen - Altersklasse B">
                  <RANKINGS>
                    <RANKING place="1" resultid="409" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6" agemax="34" agemin="18" name="Sachsen - Altersklasse A">
                  <RANKINGS>
                    <RANKING place="1" resultid="446" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7" agemax="10" agemin="7" name="offen - Altersklasse F">
                  <RANKINGS>
                    <RANKING place="1" resultid="124" />
                    <RANKING place="2" resultid="139" />
                    <RANKING place="3" resultid="273" />
                    <RANKING place="4" resultid="329" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8" agemax="11" agemin="11" name="offen - Altersklasse E">
                  <RANKINGS>
                    <RANKING place="1" resultid="143" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9" agemax="13" agemin="12" name="offen - Altersklasse D">
                  <RANKINGS>
                    <RANKING place="2" resultid="229" />
                    <RANKING place="4" resultid="233" />
                    <RANKING place="3" resultid="259" />
                    <RANKING place="5" resultid="677" />
                    <RANKING place="1" resultid="715" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10" agemax="15" agemin="14" name="offen - Altersklasse C">
                  <RANKINGS>
                    <RANKING place="2" resultid="23" />
                    <RANKING place="1" resultid="433" />
                    <RANKING place="4" resultid="673" />
                    <RANKING place="3" resultid="710" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11" agemax="17" agemin="16" name="offen - Altersklasse B">
                  <RANKINGS>
                    <RANKING place="1" resultid="409" />
                    <RANKING place="2" resultid="571" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="12" agemax="34" agemin="18" name="offen - Altersklasse A">
                  <RANKINGS>
                    <RANKING place="3" resultid="35" />
                    <RANKING place="1" resultid="446" />
                    <RANKING place="2" resultid="567" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="13" agemax="44" agemin="35" name="Sachsen - Masters AK I">
                  <RANKINGS>
                    <RANKING place="1" resultid="585" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="14" agemax="45" agemin="36" name="Sachsen - Masters AK II">
                  <RANKINGS>
                    <RANKING place="1" resultid="585" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15" agemax="55" agemin="46" name="Sachsen - Masters AK III">
                  <RANKINGS>
                    <RANKING place="1" resultid="517" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="16" agemax="65" agemin="56" name="Sachsen - Masters AK IV">
                  <RANKINGS>
                    <RANKING place="1" resultid="52" />
                    <RANKING place="2" resultid="364" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="17" agemax="-1" agemin="66" name="Sachsen - Masters AK V" />
                <AGEGROUP agegroupid="18" agemax="44" agemin="35" name="offen - Masters AK I">
                  <RANKINGS>
                    <RANKING place="1" resultid="585" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="19" agemax="45" agemin="36" name="offen - Masters AK II">
                  <RANKINGS>
                    <RANKING place="1" resultid="585" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="20" agemax="55" agemin="46" name="offen - Masters AK III">
                  <RANKINGS>
                    <RANKING place="1" resultid="517" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="21" agemax="65" agemin="56" name="offen - Masters AK IV">
                  <RANKINGS>
                    <RANKING place="1" resultid="52" />
                    <RANKING place="2" resultid="364" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="22" agemax="-1" agemin="66" name="offen - Masters AK V" />
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="3" number="3" gender="F" round="TIM">
              <SWIMSTYLE stroke="IMMERSION" technique="DIVE" relaycount="1" distance="50" />
              <FEE value="600" currency="EUR" />
              <HEATS>
                <HEAT heatid="3001" number="1" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="3" agemax="13" agemin="12" name="Sachsen - Altersklasse D">
                  <RANKINGS>
                    <RANKING place="2" resultid="287" />
                    <RANKING place="1" resultid="416" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="15" agemin="14" name="Sachsen - Altersklasse C" />
                <AGEGROUP agegroupid="9" agemax="13" agemin="12" name="offen - Altersklasse D">
                  <RANKINGS>
                    <RANKING place="1" resultid="4" />
                    <RANKING place="6" resultid="128" />
                    <RANKING place="5" resultid="287" />
                    <RANKING place="3" resultid="416" />
                    <RANKING place="2" resultid="660" />
                    <RANKING place="4" resultid="669" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10" agemax="15" agemin="14" name="offen - Altersklasse C" />
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="4" number="4" gender="M" round="TIM">
              <SWIMSTYLE stroke="IMMERSION" technique="DIVE" relaycount="1" distance="50" />
              <FEE value="600" currency="EUR" />
              <HEATS>
                <HEAT heatid="4001" number="1" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="3" agemax="13" agemin="12" name="Sachsen - Altersklasse D">
                  <RANKINGS>
                    <RANKING place="1" resultid="421" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="15" agemin="14" name="Sachsen - Altersklasse C">
                  <RANKINGS>
                    <RANKING place="1" resultid="303" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9" agemax="13" agemin="12" name="offen - Altersklasse D">
                  <RANKINGS>
                    <RANKING place="2" resultid="421" />
                    <RANKING place="1" resultid="681" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10" agemax="15" agemin="14" name="offen - Altersklasse C">
                  <RANKINGS>
                    <RANKING place="2" resultid="303" />
                    <RANKING place="1" resultid="711" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="5" number="5" gender="F" round="TIM">
              <SWIMSTYLE stroke="APNEA" relaycount="1" distance="50" />
              <FEE value="600" currency="EUR" />
              <HEATS>
                <HEAT heatid="5001" number="1" />
                <HEAT heatid="5002" number="2" />
                <HEAT heatid="5003" number="3" />
                <HEAT heatid="5004" number="4" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="4" agemax="15" agemin="14" name="Sachsen - Altersklasse C">
                  <RANKINGS>
                    <RANKING place="3" resultid="294" />
                    <RANKING place="1" resultid="333" />
                    <RANKING place="2" resultid="458" />
                    <RANKING place="4" resultid="497" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="17" agemin="16" name="Sachsen - Altersklasse B">
                  <RANKINGS>
                    <RANKING place="6" resultid="60" />
                    <RANKING place="1" resultid="297" />
                    <RANKING place="5" resultid="588" />
                    <RANKING place="2" resultid="610" />
                    <RANKING place="3" resultid="618" />
                    <RANKING place="4" resultid="630" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6" agemax="34" agemin="18" name="Sachsen - Altersklasse A">
                  <RANKINGS>
                    <RANKING place="6" resultid="338" />
                    <RANKING place="5" resultid="488" />
                    <RANKING place="3" resultid="494" />
                    <RANKING place="2" resultid="626" />
                    <RANKING place="1" resultid="639" />
                    <RANKING place="4" resultid="654" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10" agemax="15" agemin="14" name="offen - Altersklasse C">
                  <RANKINGS>
                    <RANKING place="5" resultid="31" />
                    <RANKING place="3" resultid="294" />
                    <RANKING place="1" resultid="333" />
                    <RANKING place="2" resultid="458" />
                    <RANKING place="6" resultid="497" />
                    <RANKING place="4" resultid="664" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11" agemax="17" agemin="16" name="offen - Altersklasse B">
                  <RANKINGS>
                    <RANKING place="1" resultid="13" />
                    <RANKING place="14" resultid="60" />
                    <RANKING place="3" resultid="66" />
                    <RANKING place="5" resultid="86" />
                    <RANKING place="9" resultid="237" />
                    <RANKING place="4" resultid="240" />
                    <RANKING place="8" resultid="297" />
                    <RANKING place="6" resultid="548" />
                    <RANKING place="2" resultid="562" />
                    <RANKING place="13" resultid="588" />
                    <RANKING place="10" resultid="610" />
                    <RANKING place="11" resultid="618" />
                    <RANKING place="12" resultid="630" />
                    <RANKING place="7" resultid="685" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="12" agemax="34" agemin="18" name="offen - Altersklasse A">
                  <RANKINGS>
                    <RANKING place="5" resultid="8" />
                    <RANKING place="2" resultid="69" />
                    <RANKING place="8" resultid="338" />
                    <RANKING place="7" resultid="488" />
                    <RANKING place="4" resultid="494" />
                    <RANKING place="3" resultid="626" />
                    <RANKING place="1" resultid="639" />
                    <RANKING place="6" resultid="654" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="13" agemax="44" agemin="35" name="Sachsen - Masters AK I" />
                <AGEGROUP agegroupid="14" agemax="45" agemin="36" name="Sachsen - Masters AK II" />
                <AGEGROUP agegroupid="15" agemax="55" agemin="46" name="Sachsen - Masters AK III">
                  <RANKINGS>
                    <RANKING place="1" resultid="524" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="16" agemax="65" agemin="56" name="Sachsen - Masters AK IV" />
                <AGEGROUP agegroupid="17" agemax="-1" agemin="66" name="Sachsen - Masters AK V" />
                <AGEGROUP agegroupid="18" agemax="44" agemin="35" name="offen - Masters AK I">
                  <RANKINGS>
                    <RANKING place="1" resultid="697" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="19" agemax="45" agemin="36" name="offen - Masters AK II">
                  <RANKINGS>
                    <RANKING place="1" resultid="697" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="20" agemax="55" agemin="46" name="offen - Masters AK III">
                  <RANKINGS>
                    <RANKING place="1" resultid="524" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="21" agemax="65" agemin="56" name="offen - Masters AK IV">
                  <RANKINGS>
                    <RANKING place="1" resultid="700" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="22" agemax="-1" agemin="66" name="offen - Masters AK V" />
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="6" number="6" gender="M" round="TIM">
              <SWIMSTYLE stroke="APNEA" relaycount="1" distance="50" />
              <FEE value="600" currency="EUR" />
              <HEATS>
                <HEAT heatid="6001" number="1" />
                <HEAT heatid="6002" number="2" />
                <HEAT heatid="6003" number="3" />
                <HEAT heatid="6004" number="4" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="4" agemax="15" agemin="14" name="Sachsen - Altersklasse C">
                  <RANKINGS>
                    <RANKING place="3" resultid="276" />
                    <RANKING place="2" resultid="317" />
                    <RANKING place="4" resultid="461" />
                    <RANKING place="1" resultid="481" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="17" agemin="16" name="Sachsen - Altersklasse B">
                  <RANKINGS>
                    <RANKING place="1" resultid="437" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6" agemax="34" agemin="18" name="Sachsen - Altersklasse A">
                  <RANKINGS>
                    <RANKING place="2" resultid="48" />
                    <RANKING place="1" resultid="300" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10" agemax="15" agemin="14" name="offen - Altersklasse C">
                  <RANKINGS>
                    <RANKING place="2" resultid="18" />
                    <RANKING place="4" resultid="255" />
                    <RANKING place="5" resultid="276" />
                    <RANKING place="3" resultid="317" />
                    <RANKING place="6" resultid="461" />
                    <RANKING place="1" resultid="481" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11" agemax="17" agemin="16" name="offen - Altersklasse B">
                  <RANKINGS>
                    <RANKING place="4" resultid="215" />
                    <RANKING place="2" resultid="437" />
                    <RANKING place="3" resultid="535" />
                    <RANKING place="1" resultid="689" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="12" agemax="34" agemin="18" name="offen - Altersklasse A">
                  <RANKINGS>
                    <RANKING place="4" resultid="48" />
                    <RANKING place="2" resultid="135" />
                    <RANKING place="1" resultid="300" />
                    <RANKING place="3" resultid="539" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="13" agemax="44" agemin="35" name="Sachsen - Masters AK I" />
                <AGEGROUP agegroupid="14" agemax="45" agemin="36" name="Sachsen - Masters AK II">
                  <RANKINGS>
                    <RANKING place="2" resultid="514" />
                    <RANKING place="1" resultid="598" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15" agemax="55" agemin="46" name="Sachsen - Masters AK III">
                  <RANKINGS>
                    <RANKING place="1" resultid="42" />
                    <RANKING place="2" resultid="521" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="16" agemax="65" agemin="56" name="Sachsen - Masters AK IV">
                  <RANKINGS>
                    <RANKING place="1" resultid="53" />
                    <RANKING place="2" resultid="527" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="17" agemax="-1" agemin="66" name="Sachsen - Masters AK V">
                  <RANKINGS>
                    <RANKING place="1" resultid="324" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="18" agemax="44" agemin="35" name="offen - Masters AK I" />
                <AGEGROUP agegroupid="19" agemax="45" agemin="36" name="offen - Masters AK II">
                  <RANKINGS>
                    <RANKING place="2" resultid="514" />
                    <RANKING place="1" resultid="598" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="20" agemax="55" agemin="46" name="offen - Masters AK III">
                  <RANKINGS>
                    <RANKING place="2" resultid="42" />
                    <RANKING place="3" resultid="116" />
                    <RANKING place="1" resultid="201" />
                    <RANKING place="4" resultid="521" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="21" agemax="65" agemin="56" name="offen - Masters AK IV">
                  <RANKINGS>
                    <RANKING place="1" resultid="53" />
                    <RANKING place="2" resultid="527" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="22" agemax="-1" agemin="66" name="offen - Masters AK V">
                  <RANKINGS>
                    <RANKING place="1" resultid="324" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="7" number="7" gender="F" round="TIM">
              <SWIMSTYLE stroke="SURFACE" relaycount="1" distance="100" />
              <FEE value="600" currency="EUR" />
              <HEATS>
                <HEAT heatid="7001" number="1" />
                <HEAT heatid="7002" number="2" />
                <HEAT heatid="7003" number="3" />
                <HEAT heatid="7004" number="4" />
                <HEAT heatid="7005" number="5" />
                <HEAT heatid="7006" number="6" />
                <HEAT heatid="7007" number="7" />
                <HEAT heatid="7008" number="8" />
                <HEAT heatid="7009" number="9" />
                <HEAT heatid="7010" number="10" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="10" agemin="7" name="Sachsen - Altersklasse F">
                  <RANKINGS>
                    <RANKING place="3" resultid="401" />
                    <RANKING place="2" resultid="441" />
                    <RANKING place="1" resultid="467" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2" agemax="11" agemin="11" name="Sachsen - Altersklasse E">
                  <RANKINGS>
                    <RANKING place="1" resultid="348" />
                    <RANKING place="3" resultid="379" />
                    <RANKING place="2" resultid="583" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3" agemax="13" agemin="12" name="Sachsen - Altersklasse D">
                  <RANKINGS>
                    <RANKING place="2" resultid="281" />
                    <RANKING place="7" resultid="288" />
                    <RANKING place="5" resultid="292" />
                    <RANKING place="13" resultid="341" />
                    <RANKING place="8" resultid="376" />
                    <RANKING place="6" resultid="394" />
                    <RANKING place="4" resultid="398" />
                    <RANKING place="1" resultid="417" />
                    <RANKING place="10" resultid="455" />
                    <RANKING place="15" resultid="474" />
                    <RANKING place="14" resultid="478" />
                    <RANKING place="3" resultid="491" />
                    <RANKING place="12" resultid="616" />
                    <RANKING place="11" resultid="622" />
                    <RANKING place="9" resultid="633" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="15" agemin="14" name="Sachsen - Altersklasse C">
                  <RANKINGS>
                    <RANKING place="2" resultid="334" />
                    <RANKING place="5" resultid="369" />
                    <RANKING place="3" resultid="459" />
                    <RANKING place="1" resultid="471" />
                    <RANKING place="4" resultid="498" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="17" agemin="16" name="Sachsen - Altersklasse B">
                  <RANKINGS>
                    <RANKING place="3" resultid="61" />
                    <RANKING place="5" resultid="589" />
                    <RANKING place="1" resultid="611" />
                    <RANKING place="2" resultid="619" />
                    <RANKING place="4" resultid="631" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6" agemax="34" agemin="18" name="Sachsen - Altersklasse A">
                  <RANKINGS>
                    <RANKING place="6" resultid="339" />
                    <RANKING place="5" resultid="443" />
                    <RANKING place="3" resultid="489" />
                    <RANKING place="2" resultid="495" />
                    <RANKING place="4" resultid="627" />
                    <RANKING place="1" resultid="640" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7" agemax="10" agemin="7" name="offen - Altersklasse F">
                  <RANKINGS>
                    <RANKING place="4" resultid="97" />
                    <RANKING place="6" resultid="101" />
                    <RANKING place="3" resultid="244" />
                    <RANKING place="2" resultid="247" />
                    <RANKING place="7" resultid="401" />
                    <RANKING place="5" resultid="441" />
                    <RANKING place="1" resultid="467" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8" agemax="11" agemin="11" name="offen - Altersklasse E">
                  <RANKINGS>
                    <RANKING place="1" resultid="348" />
                    <RANKING place="3" resultid="379" />
                    <RANKING place="2" resultid="583" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9" agemax="13" agemin="12" name="offen - Altersklasse D">
                  <RANKINGS>
                    <RANKING place="16" resultid="94" />
                    <RANKING place="3" resultid="281" />
                    <RANKING place="9" resultid="288" />
                    <RANKING place="6" resultid="292" />
                    <RANKING place="15" resultid="341" />
                    <RANKING place="10" resultid="376" />
                    <RANKING place="8" resultid="394" />
                    <RANKING place="5" resultid="398" />
                    <RANKING place="2" resultid="417" />
                    <RANKING place="12" resultid="455" />
                    <RANKING place="18" resultid="474" />
                    <RANKING place="17" resultid="478" />
                    <RANKING place="4" resultid="491" />
                    <RANKING place="14" resultid="616" />
                    <RANKING place="13" resultid="622" />
                    <RANKING place="11" resultid="633" />
                    <RANKING place="1" resultid="661" />
                    <RANKING place="7" resultid="670" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10" agemax="15" agemin="14" name="offen - Altersklasse C">
                  <RANKINGS>
                    <RANKING place="7" resultid="32" />
                    <RANKING place="2" resultid="334" />
                    <RANKING place="9" resultid="369" />
                    <RANKING place="5" resultid="459" />
                    <RANKING place="1" resultid="471" />
                    <RANKING place="8" resultid="498" />
                    <RANKING place="3" resultid="557" />
                    <RANKING place="4" resultid="665" />
                    <RANKING place="6" resultid="694" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11" agemax="17" agemin="16" name="offen - Altersklasse B">
                  <RANKINGS>
                    <RANKING place="2" resultid="14" />
                    <RANKING place="10" resultid="61" />
                    <RANKING place="3" resultid="67" />
                    <RANKING place="6" resultid="87" />
                    <RANKING place="4" resultid="241" />
                    <RANKING place="5" resultid="549" />
                    <RANKING place="1" resultid="563" />
                    <RANKING place="12" resultid="589" />
                    <RANKING place="8" resultid="611" />
                    <RANKING place="9" resultid="619" />
                    <RANKING place="11" resultid="631" />
                    <RANKING place="7" resultid="686" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="12" agemax="34" agemin="18" name="offen - Altersklasse A">
                  <RANKINGS>
                    <RANKING place="8" resultid="9" />
                    <RANKING place="2" resultid="70" />
                    <RANKING place="7" resultid="111" />
                    <RANKING place="10" resultid="339" />
                    <RANKING place="9" resultid="443" />
                    <RANKING place="5" resultid="489" />
                    <RANKING place="4" resultid="495" />
                    <RANKING place="3" resultid="544" />
                    <RANKING place="6" resultid="627" />
                    <RANKING place="1" resultid="640" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="13" agemax="44" agemin="35" name="Sachsen - Masters AK I">
                  <RANKINGS>
                    <RANKING place="1" resultid="509" />
                    <RANKING place="2" resultid="605" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="14" agemax="45" agemin="36" name="Sachsen - Masters AK II">
                  <RANKINGS>
                    <RANKING place="1" resultid="509" />
                    <RANKING place="2" resultid="605" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15" agemax="55" agemin="46" name="Sachsen - Masters AK III" />
                <AGEGROUP agegroupid="16" agemax="65" agemin="56" name="Sachsen - Masters AK IV">
                  <RANKINGS>
                    <RANKING place="1" resultid="357" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="17" agemax="-1" agemin="66" name="Sachsen - Masters AK V" />
                <AGEGROUP agegroupid="18" agemax="44" agemin="35" name="offen - Masters AK I">
                  <RANKINGS>
                    <RANKING place="1" resultid="509" />
                    <RANKING place="2" resultid="605" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="19" agemax="45" agemin="36" name="offen - Masters AK II">
                  <RANKINGS>
                    <RANKING place="1" resultid="509" />
                    <RANKING place="2" resultid="605" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="20" agemax="55" agemin="46" name="offen - Masters AK III">
                  <RANKINGS>
                    <RANKING place="1" resultid="198" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="21" agemax="65" agemin="56" name="offen - Masters AK IV">
                  <RANKINGS>
                    <RANKING place="2" resultid="357" />
                    <RANKING place="1" resultid="701" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="22" agemax="-1" agemin="66" name="offen - Masters AK V" />
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="8" number="8" gender="M" round="TIM">
              <SWIMSTYLE stroke="SURFACE" relaycount="1" distance="100" />
              <FEE value="600" currency="EUR" />
              <HEATS>
                <HEAT heatid="8001" number="1" />
                <HEAT heatid="8002" number="2" />
                <HEAT heatid="8003" number="3" />
                <HEAT heatid="8004" number="4" />
                <HEAT heatid="8005" number="5" />
                <HEAT heatid="8006" number="6" />
                <HEAT heatid="8007" number="7" />
                <HEAT heatid="8008" number="8" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="10" agemin="7" name="Sachsen - Altersklasse F">
                  <RANKINGS>
                    <RANKING place="2" resultid="284" />
                    <RANKING place="6" resultid="330" />
                    <RANKING place="3" resultid="351" />
                    <RANKING place="1" resultid="354" />
                    <RANKING place="4" resultid="382" />
                    <RANKING place="8" resultid="403" />
                    <RANKING place="7" resultid="407" />
                    <RANKING place="5" resultid="709" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2" agemax="11" agemin="11" name="Sachsen - Altersklasse E">
                  <RANKINGS>
                    <RANKING place="2" resultid="314" />
                    <RANKING place="1" resultid="484" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3" agemax="13" agemin="12" name="Sachsen - Altersklasse D">
                  <RANKINGS>
                    <RANKING place="1" resultid="422" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="15" agemin="14" name="Sachsen - Altersklasse C">
                  <RANKINGS>
                    <RANKING place="4" resultid="277" />
                    <RANKING place="8" resultid="304" />
                    <RANKING place="3" resultid="318" />
                    <RANKING place="2" resultid="434" />
                    <RANKING place="5" resultid="462" />
                    <RANKING place="1" resultid="482" />
                    <RANKING place="7" resultid="602" />
                    <RANKING place="6" resultid="608" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="17" agemin="16" name="Sachsen - Altersklasse B">
                  <RANKINGS>
                    <RANKING place="3" resultid="40" />
                    <RANKING place="1" resultid="410" />
                    <RANKING place="2" resultid="438" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6" agemax="34" agemin="18" name="Sachsen - Altersklasse A">
                  <RANKINGS>
                    <RANKING place="1" resultid="49" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7" agemax="10" agemin="7" name="offen - Altersklasse F">
                  <RANKINGS>
                    <RANKING place="13" resultid="114" />
                    <RANKING place="3" resultid="125" />
                    <RANKING place="10" resultid="132" />
                    <RANKING place="4" resultid="140" />
                    <RANKING place="2" resultid="226" />
                    <RANKING place="5" resultid="284" />
                    <RANKING place="9" resultid="330" />
                    <RANKING place="6" resultid="351" />
                    <RANKING place="1" resultid="354" />
                    <RANKING place="7" resultid="382" />
                    <RANKING place="12" resultid="403" />
                    <RANKING place="11" resultid="407" />
                    <RANKING place="8" resultid="709" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8" agemax="11" agemin="11" name="offen - Altersklasse E">
                  <RANKINGS>
                    <RANKING place="2" resultid="144" />
                    <RANKING place="3" resultid="263" />
                    <RANKING place="4" resultid="314" />
                    <RANKING place="1" resultid="484" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9" agemax="13" agemin="12" name="offen - Altersklasse D">
                  <RANKINGS>
                    <RANKING place="4" resultid="230" />
                    <RANKING place="5" resultid="234" />
                    <RANKING place="6" resultid="260" />
                    <RANKING place="3" resultid="422" />
                    <RANKING place="7" resultid="678" />
                    <RANKING place="2" resultid="682" />
                    <RANKING place="1" resultid="716" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10" agemax="15" agemin="14" name="offen - Altersklasse C">
                  <RANKINGS>
                    <RANKING place="5" resultid="19" />
                    <RANKING place="3" resultid="256" />
                    <RANKING place="7" resultid="277" />
                    <RANKING place="12" resultid="304" />
                    <RANKING place="4" resultid="318" />
                    <RANKING place="2" resultid="434" />
                    <RANKING place="9" resultid="462" />
                    <RANKING place="1" resultid="482" />
                    <RANKING place="11" resultid="602" />
                    <RANKING place="10" resultid="608" />
                    <RANKING place="6" resultid="674" />
                    <RANKING place="8" resultid="712" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11" agemax="17" agemin="16" name="offen - Altersklasse B">
                  <RANKINGS>
                    <RANKING place="5" resultid="40" />
                    <RANKING place="2" resultid="410" />
                    <RANKING place="3" resultid="438" />
                    <RANKING place="4" resultid="536" />
                    <RANKING place="1" resultid="690" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="12" agemax="34" agemin="18" name="offen - Altersklasse A">
                  <RANKINGS>
                    <RANKING place="4" resultid="49" />
                    <RANKING place="2" resultid="136" />
                    <RANKING place="1" resultid="540" />
                    <RANKING place="3" resultid="568" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="13" agemax="44" agemin="35" name="Sachsen - Masters AK I">
                  <RANKINGS>
                    <RANKING place="1" resultid="586" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="14" agemax="45" agemin="36" name="Sachsen - Masters AK II">
                  <RANKINGS>
                    <RANKING place="2" resultid="515" />
                    <RANKING place="1" resultid="586" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15" agemax="55" agemin="46" name="Sachsen - Masters AK III">
                  <RANKINGS>
                    <RANKING place="2" resultid="43" />
                    <RANKING place="1" resultid="518" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="16" agemax="65" agemin="56" name="Sachsen - Masters AK IV">
                  <RANKINGS>
                    <RANKING place="1" resultid="54" />
                    <RANKING place="3" resultid="365" />
                    <RANKING place="2" resultid="528" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="17" agemax="-1" agemin="66" name="Sachsen - Masters AK V">
                  <RANKINGS>
                    <RANKING place="1" resultid="325" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="18" agemax="44" agemin="35" name="offen - Masters AK I">
                  <RANKINGS>
                    <RANKING place="1" resultid="586" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="19" agemax="45" agemin="36" name="offen - Masters AK II">
                  <RANKINGS>
                    <RANKING place="2" resultid="515" />
                    <RANKING place="1" resultid="586" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="20" agemax="55" agemin="46" name="offen - Masters AK III">
                  <RANKINGS>
                    <RANKING place="3" resultid="43" />
                    <RANKING place="4" resultid="117" />
                    <RANKING place="2" resultid="202" />
                    <RANKING place="1" resultid="518" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="21" agemax="65" agemin="56" name="offen - Masters AK IV">
                  <RANKINGS>
                    <RANKING place="1" resultid="54" />
                    <RANKING place="3" resultid="365" />
                    <RANKING place="2" resultid="528" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="22" agemax="-1" agemin="66" name="offen - Masters AK V">
                  <RANKINGS>
                    <RANKING place="1" resultid="325" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="9" number="9" gender="F" round="TIM">
              <SWIMSTYLE stroke="SURFACE" relaycount="1" distance="800" />
              <FEE value="600" currency="EUR" />
              <HEATS>
                <HEAT heatid="9001" number="1" />
                <HEAT heatid="9002" number="2" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="2" agemax="11" agemin="11" name="Sachsen - Altersklasse E" />
                <AGEGROUP agegroupid="3" agemax="13" agemin="12" name="Sachsen - Altersklasse D" />
                <AGEGROUP agegroupid="4" agemax="15" agemin="14" name="Sachsen - Altersklasse C">
                  <RANKINGS>
                    <RANKING place="1" resultid="707" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="17" agemin="16" name="Sachsen - Altersklasse B">
                  <RANKINGS>
                    <RANKING place="1" resultid="298" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6" agemax="34" agemin="18" name="Sachsen - Altersklasse A">
                  <RANKINGS>
                    <RANKING place="2" resultid="414" />
                    <RANKING place="1" resultid="721" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8" agemax="11" agemin="11" name="offen - Altersklasse E" />
                <AGEGROUP agegroupid="9" agemax="13" agemin="12" name="offen - Altersklasse D">
                  <RANKINGS>
                    <RANKING place="1" resultid="5" />
                    <RANKING place="2" resultid="129" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10" agemax="15" agemin="14" name="offen - Altersklasse C">
                  <RANKINGS>
                    <RANKING place="1" resultid="558" />
                    <RANKING place="2" resultid="707" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11" agemax="17" agemin="16" name="offen - Altersklasse B">
                  <RANKINGS>
                    <RANKING place="2" resultid="252" />
                    <RANKING place="3" resultid="298" />
                    <RANKING place="1" resultid="564" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="12" agemax="34" agemin="18" name="offen - Altersklasse A">
                  <RANKINGS>
                    <RANKING place="2" resultid="28" />
                    <RANKING place="3" resultid="414" />
                    <RANKING place="1" resultid="721" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="13" agemax="44" agemin="35" name="Sachsen - Masters AK I" />
                <AGEGROUP agegroupid="14" agemax="45" agemin="36" name="Sachsen - Masters AK II" />
                <AGEGROUP agegroupid="15" agemax="55" agemin="46" name="Sachsen - Masters AK III" />
                <AGEGROUP agegroupid="16" agemax="65" agemin="56" name="Sachsen - Masters AK IV" />
                <AGEGROUP agegroupid="17" agemax="-1" agemin="66" name="Sachsen - Masters AK V" />
                <AGEGROUP agegroupid="18" agemax="44" agemin="35" name="offen - Masters AK I" />
                <AGEGROUP agegroupid="19" agemax="45" agemin="36" name="offen - Masters AK II" />
                <AGEGROUP agegroupid="20" agemax="55" agemin="46" name="offen - Masters AK III" />
                <AGEGROUP agegroupid="21" agemax="65" agemin="56" name="offen - Masters AK IV" />
                <AGEGROUP agegroupid="22" agemax="-1" agemin="66" name="offen - Masters AK V" />
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="10" number="10" gender="M" round="TIM">
              <SWIMSTYLE stroke="SURFACE" relaycount="1" distance="800" />
              <FEE value="600" currency="EUR" />
              <HEATS>
                <HEAT heatid="10000" number="0" />
                <HEAT heatid="10001" number="1" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="2" agemax="11" agemin="11" name="Sachsen - Altersklasse E" />
                <AGEGROUP agegroupid="3" agemax="13" agemin="12" name="Sachsen - Altersklasse D" />
                <AGEGROUP agegroupid="4" agemax="15" agemin="14" name="Sachsen - Altersklasse C" />
                <AGEGROUP agegroupid="5" agemax="17" agemin="16" name="Sachsen - Altersklasse B" />
                <AGEGROUP agegroupid="6" agemax="34" agemin="18" name="Sachsen - Altersklasse A">
                  <RANKINGS>
                    <RANKING place="1" resultid="447" />
                    <RANKING place="2" resultid="452" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8" agemax="11" agemin="11" name="offen - Altersklasse E" />
                <AGEGROUP agegroupid="9" agemax="13" agemin="12" name="offen - Altersklasse D" />
                <AGEGROUP agegroupid="10" agemax="15" agemin="14" name="offen - Altersklasse C">
                  <RANKINGS>
                    <RANKING place="1" resultid="20" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11" agemax="17" agemin="16" name="offen - Altersklasse B">
                  <RANKINGS>
                    <RANKING place="1" resultid="572" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="12" agemax="34" agemin="18" name="offen - Altersklasse A">
                  <RANKINGS>
                    <RANKING place="2" resultid="1" />
                    <RANKING place="4" resultid="36" />
                    <RANKING place="1" resultid="447" />
                    <RANKING place="3" resultid="452" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="13" agemax="44" agemin="35" name="Sachsen - Masters AK I" />
                <AGEGROUP agegroupid="14" agemax="45" agemin="36" name="Sachsen - Masters AK II" />
                <AGEGROUP agegroupid="15" agemax="55" agemin="46" name="Sachsen - Masters AK III" />
                <AGEGROUP agegroupid="16" agemax="65" agemin="56" name="Sachsen - Masters AK IV">
                  <RANKINGS>
                    <RANKING place="1" resultid="55" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="17" agemax="-1" agemin="66" name="Sachsen - Masters AK V" />
                <AGEGROUP agegroupid="18" agemax="44" agemin="35" name="offen - Masters AK I" />
                <AGEGROUP agegroupid="19" agemax="45" agemin="36" name="offen - Masters AK II" />
                <AGEGROUP agegroupid="20" agemax="55" agemin="46" name="offen - Masters AK III" />
                <AGEGROUP agegroupid="21" agemax="65" agemin="56" name="offen - Masters AK IV">
                  <RANKINGS>
                    <RANKING place="1" resultid="55" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="22" agemax="-1" agemin="66" name="offen - Masters AK V" />
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="11" number="11" gender="F" round="TIM">
              <SWIMSTYLE stroke="BIFIN" relaycount="1" distance="50" />
              <FEE value="600" currency="EUR" />
              <HEATS>
                <HEAT heatid="11001" number="1" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="13" agemax="44" agemin="35" name="Sachsen - Masters AK I">
                  <RANKINGS>
                    <RANKING place="1" resultid="510" />
                    <RANKING place="2" resultid="512" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="14" agemax="45" agemin="36" name="Sachsen - Masters AK II">
                  <RANKINGS>
                    <RANKING place="1" resultid="510" />
                    <RANKING place="2" resultid="512" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15" agemax="55" agemin="46" name="Sachsen - Masters AK III">
                  <RANKINGS>
                    <RANKING place="1" resultid="505" />
                    <RANKING place="2" resultid="525" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="16" agemax="65" agemin="56" name="Sachsen - Masters AK IV">
                  <RANKINGS>
                    <RANKING place="1" resultid="507" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="17" agemax="-1" agemin="66" name="Sachsen - Masters AK V" />
                <AGEGROUP agegroupid="18" agemax="44" agemin="35" name="offen - Masters AK I">
                  <RANKINGS>
                    <RANKING place="1" resultid="510" />
                    <RANKING place="2" resultid="512" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="19" agemax="45" agemin="36" name="offen - Masters AK II">
                  <RANKINGS>
                    <RANKING place="1" resultid="510" />
                    <RANKING place="2" resultid="512" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="20" agemax="55" agemin="46" name="offen - Masters AK III">
                  <RANKINGS>
                    <RANKING place="1" resultid="505" />
                    <RANKING place="2" resultid="525" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="21" agemax="65" agemin="56" name="offen - Masters AK IV">
                  <RANKINGS>
                    <RANKING place="2" resultid="507" />
                    <RANKING place="1" resultid="702" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="22" agemax="-1" agemin="66" name="offen - Masters AK V" />
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="12" number="12" gender="M" round="TIM">
              <SWIMSTYLE stroke="BIFIN" relaycount="1" distance="50" />
              <FEE value="600" currency="EUR" />
              <HEATS>
                <HEAT heatid="12001" number="1" />
                <HEAT heatid="12002" number="2" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="13" agemax="44" agemin="35" name="Sachsen - Masters AK I" />
                <AGEGROUP agegroupid="14" agemax="45" agemin="36" name="Sachsen - Masters AK II">
                  <RANKINGS>
                    <RANKING place="2" resultid="516" />
                    <RANKING place="1" resultid="599" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15" agemax="55" agemin="46" name="Sachsen - Masters AK III">
                  <RANKINGS>
                    <RANKING place="2" resultid="64" />
                    <RANKING place="1" resultid="372" />
                    <RANKING place="3" resultid="522" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="16" agemax="65" agemin="56" name="Sachsen - Masters AK IV">
                  <RANKINGS>
                    <RANKING place="2" resultid="366" />
                    <RANKING place="1" resultid="529" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="17" agemax="-1" agemin="66" name="Sachsen - Masters AK V">
                  <RANKINGS>
                    <RANKING place="1" resultid="326" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="18" agemax="44" agemin="35" name="offen - Masters AK I" />
                <AGEGROUP agegroupid="19" agemax="45" agemin="36" name="offen - Masters AK II">
                  <RANKINGS>
                    <RANKING place="2" resultid="516" />
                    <RANKING place="1" resultid="599" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="20" agemax="55" agemin="46" name="offen - Masters AK III">
                  <RANKINGS>
                    <RANKING place="2" resultid="64" />
                    <RANKING place="3" resultid="203" />
                    <RANKING place="1" resultid="372" />
                    <RANKING place="4" resultid="522" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="21" agemax="65" agemin="56" name="offen - Masters AK IV">
                  <RANKINGS>
                    <RANKING place="2" resultid="366" />
                    <RANKING place="1" resultid="529" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="22" agemax="-1" agemin="66" name="offen - Masters AK V">
                  <RANKINGS>
                    <RANKING place="1" resultid="326" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="13" number="13" gender="X" round="TIM">
              <SWIMSTYLE stroke="SURFACE" relaycount="4" distance="50" />
              <FEE value="800" currency="EUR" />
              <HEATS>
                <HEAT heatid="13001" number="1" />
                <HEAT heatid="13002" number="2" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="3" agemax="-1" agemin="7" name="Sachsen - offene Wertung">
                  <RANKINGS>
                    <RANKING place="2" resultid="269" />
                    <RANKING place="7" resultid="272" />
                    <RANKING place="5" resultid="321" />
                    <RANKING place="8" resultid="323" />
                    <RANKING place="1" resultid="426" />
                    <RANKING place="6" resultid="430" />
                    <RANKING place="9" resultid="432" />
                    <RANKING place="3" resultid="504" />
                    <RANKING place="4" resultid="582" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6" agemax="-1" agemin="7" name="offen - offene Wertung">
                  <RANKINGS>
                    <RANKING place="4" resultid="266" />
                    <RANKING place="12" resultid="267" />
                    <RANKING place="3" resultid="269" />
                    <RANKING place="10" resultid="272" />
                    <RANKING place="8" resultid="321" />
                    <RANKING place="11" resultid="323" />
                    <RANKING place="2" resultid="426" />
                    <RANKING place="9" resultid="430" />
                    <RANKING place="13" resultid="432" />
                    <RANKING place="5" resultid="504" />
                    <RANKING place="7" resultid="582" />
                    <RANKING place="6" resultid="658" />
                    <RANKING place="1" resultid="720" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
          </EVENTS>
        </SESSION>
        <SESSION number="2" date="2023-04-01" daytime="00:52">
          <EVENTS>
            <EVENT eventid="14" number="14" gender="F" round="TIM">
              <SWIMSTYLE stroke="SURFACE" relaycount="1" distance="50" />
              <FEE value="600" currency="EUR" />
              <HEATS>
                <HEAT heatid="14001" number="1" />
                <HEAT heatid="14002" number="2" />
                <HEAT heatid="14003" number="3" />
                <HEAT heatid="14004" number="4" />
                <HEAT heatid="14005" number="5" />
                <HEAT heatid="14006" number="6" />
                <HEAT heatid="14007" number="7" />
                <HEAT heatid="14008" number="8" />
                <HEAT heatid="14009" number="9" />
                <HEAT heatid="14010" number="10" />
                <HEAT heatid="14011" number="11" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="10" agemin="7" name="Sachsen - Altersklasse F">
                  <RANKINGS>
                    <RANKING place="5" resultid="402" />
                    <RANKING place="4" resultid="442" />
                    <RANKING place="3" resultid="468" />
                    <RANKING place="1" resultid="501" />
                    <RANKING place="2" resultid="649" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2" agemax="11" agemin="11" name="Sachsen - Altersklasse E">
                  <RANKINGS>
                    <RANKING place="1" resultid="349" />
                    <RANKING place="3" resultid="380" />
                    <RANKING place="2" resultid="584" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3" agemax="13" agemin="12" name="Sachsen - Altersklasse D">
                  <RANKINGS>
                    <RANKING place="2" resultid="282" />
                    <RANKING place="7" resultid="289" />
                    <RANKING place="14" resultid="342" />
                    <RANKING place="6" resultid="377" />
                    <RANKING place="4" resultid="399" />
                    <RANKING place="3" resultid="418" />
                    <RANKING place="8" resultid="456" />
                    <RANKING place="13" resultid="475" />
                    <RANKING place="12" resultid="479" />
                    <RANKING place="1" resultid="492" />
                    <RANKING place="11" resultid="615" />
                    <RANKING place="9" resultid="617" />
                    <RANKING place="10" resultid="623" />
                    <RANKING place="5" resultid="634" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="15" agemin="14" name="Sachsen - Altersklasse C">
                  <RANKINGS>
                    <RANKING place="3" resultid="295" />
                    <RANKING place="2" resultid="335" />
                    <RANKING place="5" resultid="370" />
                    <RANKING place="1" resultid="472" />
                    <RANKING place="4" resultid="499" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="17" agemin="16" name="Sachsen - Altersklasse B">
                  <RANKINGS>
                    <RANKING place="4" resultid="62" />
                    <RANKING place="1" resultid="465" />
                    <RANKING place="6" resultid="590" />
                    <RANKING place="2" resultid="612" />
                    <RANKING place="3" resultid="620" />
                    <RANKING place="5" resultid="632" />
                    <RANKING place="7" resultid="644" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6" agemax="34" agemin="18" name="Sachsen - Altersklasse A">
                  <RANKINGS>
                    <RANKING place="5" resultid="340" />
                    <RANKING place="3" resultid="444" />
                    <RANKING place="4" resultid="496" />
                    <RANKING place="2" resultid="628" />
                    <RANKING place="1" resultid="641" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7" agemax="10" agemin="7" name="offen - Altersklasse F">
                  <RANKINGS>
                    <RANKING place="7" resultid="98" />
                    <RANKING place="6" resultid="102" />
                    <RANKING place="5" resultid="245" />
                    <RANKING place="4" resultid="248" />
                    <RANKING place="9" resultid="402" />
                    <RANKING place="8" resultid="442" />
                    <RANKING place="3" resultid="468" />
                    <RANKING place="1" resultid="501" />
                    <RANKING place="2" resultid="649" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8" agemax="11" agemin="11" name="offen - Altersklasse E">
                  <RANKINGS>
                    <RANKING place="1" resultid="349" />
                    <RANKING place="3" resultid="380" />
                    <RANKING place="2" resultid="584" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9" agemax="13" agemin="12" name="offen - Altersklasse D">
                  <RANKINGS>
                    <RANKING place="1" resultid="6" />
                    <RANKING place="19" resultid="95" />
                    <RANKING place="13" resultid="130" />
                    <RANKING place="4" resultid="282" />
                    <RANKING place="10" resultid="289" />
                    <RANKING place="18" resultid="342" />
                    <RANKING place="9" resultid="377" />
                    <RANKING place="6" resultid="399" />
                    <RANKING place="5" resultid="418" />
                    <RANKING place="11" resultid="456" />
                    <RANKING place="17" resultid="475" />
                    <RANKING place="16" resultid="479" />
                    <RANKING place="3" resultid="492" />
                    <RANKING place="15" resultid="615" />
                    <RANKING place="12" resultid="617" />
                    <RANKING place="14" resultid="623" />
                    <RANKING place="7" resultid="634" />
                    <RANKING place="2" resultid="662" />
                    <RANKING place="8" resultid="671" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10" agemax="15" agemin="14" name="offen - Altersklasse C">
                  <RANKINGS>
                    <RANKING place="4" resultid="295" />
                    <RANKING place="3" resultid="335" />
                    <RANKING place="8" resultid="370" />
                    <RANKING place="1" resultid="472" />
                    <RANKING place="7" resultid="499" />
                    <RANKING place="2" resultid="559" />
                    <RANKING place="5" resultid="666" />
                    <RANKING place="6" resultid="695" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11" agemax="17" agemin="16" name="offen - Altersklasse B">
                  <RANKINGS>
                    <RANKING place="2" resultid="15" />
                    <RANKING place="13" resultid="62" />
                    <RANKING place="6" resultid="88" />
                    <RANKING place="1" resultid="147" />
                    <RANKING place="10" resultid="239" />
                    <RANKING place="5" resultid="242" />
                    <RANKING place="8" resultid="253" />
                    <RANKING place="7" resultid="465" />
                    <RANKING place="4" resultid="550" />
                    <RANKING place="3" resultid="565" />
                    <RANKING place="15" resultid="590" />
                    <RANKING place="11" resultid="612" />
                    <RANKING place="12" resultid="620" />
                    <RANKING place="14" resultid="632" />
                    <RANKING place="16" resultid="644" />
                    <RANKING place="9" resultid="687" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="12" agemax="34" agemin="18" name="offen - Altersklasse A">
                  <RANKINGS>
                    <RANKING place="2" resultid="71" />
                    <RANKING place="4" resultid="112" />
                    <RANKING place="8" resultid="340" />
                    <RANKING place="6" resultid="444" />
                    <RANKING place="7" resultid="496" />
                    <RANKING place="5" resultid="545" />
                    <RANKING place="3" resultid="628" />
                    <RANKING place="1" resultid="641" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="13" agemax="44" agemin="35" name="Sachsen - Masters AK I">
                  <RANKINGS>
                    <RANKING place="1" resultid="511" />
                    <RANKING place="3" resultid="513" />
                    <RANKING place="2" resultid="606" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="14" agemax="45" agemin="36" name="Sachsen - Masters AK II">
                  <RANKINGS>
                    <RANKING place="1" resultid="511" />
                    <RANKING place="3" resultid="513" />
                    <RANKING place="2" resultid="606" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15" agemax="55" agemin="46" name="Sachsen - Masters AK III">
                  <RANKINGS>
                    <RANKING place="2" resultid="506" />
                    <RANKING place="1" resultid="526" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="16" agemax="65" agemin="56" name="Sachsen - Masters AK IV">
                  <RANKINGS>
                    <RANKING place="2" resultid="358" />
                    <RANKING place="1" resultid="508" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="17" agemax="-1" agemin="66" name="Sachsen - Masters AK V">
                  <RANKINGS>
                    <RANKING place="1" resultid="362" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="18" agemax="44" agemin="35" name="offen - Masters AK I">
                  <RANKINGS>
                    <RANKING place="1" resultid="511" />
                    <RANKING place="4" resultid="513" />
                    <RANKING place="3" resultid="606" />
                    <RANKING place="2" resultid="698" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="19" agemax="45" agemin="36" name="offen - Masters AK II">
                  <RANKINGS>
                    <RANKING place="1" resultid="511" />
                    <RANKING place="4" resultid="513" />
                    <RANKING place="3" resultid="606" />
                    <RANKING place="2" resultid="698" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="20" agemax="55" agemin="46" name="offen - Masters AK III">
                  <RANKINGS>
                    <RANKING place="2" resultid="199" />
                    <RANKING place="3" resultid="506" />
                    <RANKING place="1" resultid="526" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="21" agemax="65" agemin="56" name="offen - Masters AK IV">
                  <RANKINGS>
                    <RANKING place="3" resultid="358" />
                    <RANKING place="1" resultid="508" />
                    <RANKING place="2" resultid="703" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="22" agemax="-1" agemin="66" name="offen - Masters AK V">
                  <RANKINGS>
                    <RANKING place="1" resultid="362" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="15" number="15" gender="M" round="TIM">
              <SWIMSTYLE stroke="SURFACE" relaycount="1" distance="50" />
              <FEE value="600" currency="EUR" />
              <HEATS>
                <HEAT heatid="15001" number="1" />
                <HEAT heatid="15002" number="2" />
                <HEAT heatid="15003" number="3" />
                <HEAT heatid="15004" number="4" />
                <HEAT heatid="15005" number="5" />
                <HEAT heatid="15006" number="6" />
                <HEAT heatid="15007" number="7" />
                <HEAT heatid="15008" number="8" />
                <HEAT heatid="15009" number="9" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="10" agemin="7" name="Sachsen - Altersklasse F">
                  <RANKINGS>
                    <RANKING place="1" resultid="274" />
                    <RANKING place="3" resultid="285" />
                    <RANKING place="7" resultid="331" />
                    <RANKING place="4" resultid="352" />
                    <RANKING place="2" resultid="355" />
                    <RANKING place="5" resultid="383" />
                    <RANKING place="9" resultid="404" />
                    <RANKING place="8" resultid="408" />
                    <RANKING place="6" resultid="436" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2" agemax="11" agemin="11" name="Sachsen - Altersklasse E">
                  <RANKINGS>
                    <RANKING place="2" resultid="315" />
                    <RANKING place="1" resultid="485" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3" agemax="13" agemin="12" name="Sachsen - Altersklasse D">
                  <RANKINGS>
                    <RANKING place="1" resultid="423" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="15" agemin="14" name="Sachsen - Altersklasse C">
                  <RANKINGS>
                    <RANKING place="3" resultid="278" />
                    <RANKING place="7" resultid="305" />
                    <RANKING place="2" resultid="319" />
                    <RANKING place="4" resultid="463" />
                    <RANKING place="1" resultid="483" />
                    <RANKING place="5" resultid="603" />
                    <RANKING place="6" resultid="609" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="17" agemin="16" name="Sachsen - Altersklasse B">
                  <RANKINGS>
                    <RANKING place="3" resultid="41" />
                    <RANKING place="1" resultid="411" />
                    <RANKING place="2" resultid="439" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6" agemax="34" agemin="18" name="Sachsen - Altersklasse A">
                  <RANKINGS>
                    <RANKING place="3" resultid="50" />
                    <RANKING place="1" resultid="301" />
                    <RANKING place="2" resultid="453" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7" agemax="10" agemin="7" name="offen - Altersklasse F">
                  <RANKINGS>
                    <RANKING place="1" resultid="126" />
                    <RANKING place="10" resultid="133" />
                    <RANKING place="3" resultid="141" />
                    <RANKING place="4" resultid="227" />
                    <RANKING place="2" resultid="274" />
                    <RANKING place="6" resultid="285" />
                    <RANKING place="11" resultid="331" />
                    <RANKING place="7" resultid="352" />
                    <RANKING place="5" resultid="355" />
                    <RANKING place="8" resultid="383" />
                    <RANKING place="13" resultid="404" />
                    <RANKING place="12" resultid="408" />
                    <RANKING place="9" resultid="436" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8" agemax="11" agemin="11" name="offen - Altersklasse E">
                  <RANKINGS>
                    <RANKING place="2" resultid="145" />
                    <RANKING place="3" resultid="264" />
                    <RANKING place="4" resultid="315" />
                    <RANKING place="1" resultid="485" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9" agemax="13" agemin="12" name="offen - Altersklasse D">
                  <RANKINGS>
                    <RANKING place="8" resultid="220" />
                    <RANKING place="4" resultid="231" />
                    <RANKING place="5" resultid="235" />
                    <RANKING place="6" resultid="261" />
                    <RANKING place="3" resultid="423" />
                    <RANKING place="7" resultid="679" />
                    <RANKING place="2" resultid="683" />
                    <RANKING place="1" resultid="717" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10" agemax="15" agemin="14" name="offen - Altersklasse C">
                  <RANKINGS>
                    <RANKING place="2" resultid="257" />
                    <RANKING place="5" resultid="278" />
                    <RANKING place="10" resultid="305" />
                    <RANKING place="3" resultid="319" />
                    <RANKING place="7" resultid="463" />
                    <RANKING place="1" resultid="483" />
                    <RANKING place="8" resultid="603" />
                    <RANKING place="9" resultid="609" />
                    <RANKING place="6" resultid="675" />
                    <RANKING place="4" resultid="713" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11" agemax="17" agemin="16" name="offen - Altersklasse B">
                  <RANKINGS>
                    <RANKING place="6" resultid="41" />
                    <RANKING place="2" resultid="411" />
                    <RANKING place="3" resultid="439" />
                    <RANKING place="4" resultid="537" />
                    <RANKING place="5" resultid="573" />
                    <RANKING place="1" resultid="691" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="12" agemax="34" agemin="18" name="offen - Altersklasse A">
                  <RANKINGS>
                    <RANKING place="6" resultid="50" />
                    <RANKING place="4" resultid="137" />
                    <RANKING place="1" resultid="301" />
                    <RANKING place="2" resultid="453" />
                    <RANKING place="5" resultid="569" />
                    <RANKING place="3" resultid="651" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="13" agemax="44" agemin="35" name="Sachsen - Masters AK I" />
                <AGEGROUP agegroupid="14" agemax="45" agemin="36" name="Sachsen - Masters AK II">
                  <RANKINGS>
                    <RANKING place="1" resultid="600" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15" agemax="55" agemin="46" name="Sachsen - Masters AK III">
                  <RANKINGS>
                    <RANKING place="3" resultid="45" />
                    <RANKING place="2" resultid="373" />
                    <RANKING place="1" resultid="519" />
                    <RANKING place="4" resultid="523" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="16" agemax="65" agemin="56" name="Sachsen - Masters AK IV">
                  <RANKINGS>
                    <RANKING place="2" resultid="56" />
                    <RANKING place="3" resultid="367" />
                    <RANKING place="1" resultid="530" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="17" agemax="-1" agemin="66" name="Sachsen - Masters AK V">
                  <RANKINGS>
                    <RANKING place="1" resultid="327" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="18" agemax="44" agemin="35" name="offen - Masters AK I" />
                <AGEGROUP agegroupid="19" agemax="45" agemin="36" name="offen - Masters AK II">
                  <RANKINGS>
                    <RANKING place="1" resultid="600" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="20" agemax="55" agemin="46" name="offen - Masters AK III">
                  <RANKINGS>
                    <RANKING place="4" resultid="45" />
                    <RANKING place="6" resultid="118" />
                    <RANKING place="3" resultid="204" />
                    <RANKING place="2" resultid="373" />
                    <RANKING place="1" resultid="519" />
                    <RANKING place="5" resultid="523" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="21" agemax="65" agemin="56" name="offen - Masters AK IV">
                  <RANKINGS>
                    <RANKING place="2" resultid="56" />
                    <RANKING place="3" resultid="367" />
                    <RANKING place="1" resultid="530" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="22" agemax="-1" agemin="66" name="offen - Masters AK V">
                  <RANKINGS>
                    <RANKING place="1" resultid="327" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="16" number="16" gender="F" round="TIM">
              <SWIMSTYLE stroke="SURFACE" relaycount="1" distance="1500" />
              <FEE value="600" currency="EUR" />
              <HEATS>
                <HEAT heatid="16001" number="1" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="2" agemax="11" agemin="11" name="Sachsen - Altersklasse E" />
                <AGEGROUP agegroupid="3" agemax="13" agemin="12" name="Sachsen - Altersklasse D" />
                <AGEGROUP agegroupid="4" agemax="15" agemin="14" name="Sachsen - Altersklasse C" />
                <AGEGROUP agegroupid="5" agemax="17" agemin="16" name="Sachsen - Altersklasse B" />
                <AGEGROUP agegroupid="6" agemax="34" agemin="18" name="Sachsen - Altersklasse A" />
                <AGEGROUP agegroupid="8" agemax="11" agemin="11" name="offen - Altersklasse E" />
                <AGEGROUP agegroupid="9" agemax="13" agemin="12" name="offen - Altersklasse D" />
                <AGEGROUP agegroupid="10" agemax="15" agemin="14" name="offen - Altersklasse C" />
                <AGEGROUP agegroupid="11" agemax="17" agemin="16" name="offen - Altersklasse B" />
                <AGEGROUP agegroupid="12" agemax="34" agemin="18" name="offen - Altersklasse A">
                  <RANKINGS>
                    <RANKING place="1" resultid="29" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="13" agemax="44" agemin="35" name="Sachsen - Masters AK I" />
                <AGEGROUP agegroupid="14" agemax="45" agemin="36" name="Sachsen - Masters AK II" />
                <AGEGROUP agegroupid="15" agemax="55" agemin="46" name="Sachsen - Masters AK III" />
                <AGEGROUP agegroupid="16" agemax="65" agemin="56" name="Sachsen - Masters AK IV" />
                <AGEGROUP agegroupid="17" agemax="-1" agemin="66" name="Sachsen - Masters AK V" />
                <AGEGROUP agegroupid="18" agemax="44" agemin="35" name="offen - Masters AK I" />
                <AGEGROUP agegroupid="19" agemax="45" agemin="36" name="offen - Masters AK II" />
                <AGEGROUP agegroupid="20" agemax="55" agemin="46" name="offen - Masters AK III" />
                <AGEGROUP agegroupid="21" agemax="65" agemin="56" name="offen - Masters AK IV" />
                <AGEGROUP agegroupid="22" agemax="-1" agemin="66" name="offen - Masters AK V" />
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="17" number="17" gender="M" round="TIM">
              <SWIMSTYLE stroke="SURFACE" relaycount="1" distance="1500" />
              <FEE value="600" currency="EUR" />
              <HEATS>
                <HEAT heatid="17001" number="1" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="2" agemax="11" agemin="11" name="Sachsen - Altersklasse E" />
                <AGEGROUP agegroupid="3" agemax="13" agemin="12" name="Sachsen - Altersklasse D" />
                <AGEGROUP agegroupid="4" agemax="15" agemin="14" name="Sachsen - Altersklasse C" />
                <AGEGROUP agegroupid="5" agemax="17" agemin="16" name="Sachsen - Altersklasse B" />
                <AGEGROUP agegroupid="6" agemax="34" agemin="18" name="Sachsen - Altersklasse A" />
                <AGEGROUP agegroupid="8" agemax="11" agemin="11" name="offen - Altersklasse E" />
                <AGEGROUP agegroupid="9" agemax="13" agemin="12" name="offen - Altersklasse D" />
                <AGEGROUP agegroupid="10" agemax="15" agemin="14" name="offen - Altersklasse C" />
                <AGEGROUP agegroupid="11" agemax="17" agemin="16" name="offen - Altersklasse B" />
                <AGEGROUP agegroupid="12" agemax="34" agemin="18" name="offen - Altersklasse A">
                  <RANKINGS>
                    <RANKING place="1" resultid="2" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="13" agemax="44" agemin="35" name="Sachsen - Masters AK I" />
                <AGEGROUP agegroupid="14" agemax="45" agemin="36" name="Sachsen - Masters AK II" />
                <AGEGROUP agegroupid="15" agemax="55" agemin="46" name="Sachsen - Masters AK III" />
                <AGEGROUP agegroupid="16" agemax="65" agemin="56" name="Sachsen - Masters AK IV" />
                <AGEGROUP agegroupid="17" agemax="-1" agemin="66" name="Sachsen - Masters AK V" />
                <AGEGROUP agegroupid="18" agemax="44" agemin="35" name="offen - Masters AK I" />
                <AGEGROUP agegroupid="19" agemax="45" agemin="36" name="offen - Masters AK II" />
                <AGEGROUP agegroupid="20" agemax="55" agemin="46" name="offen - Masters AK III" />
                <AGEGROUP agegroupid="21" agemax="65" agemin="56" name="offen - Masters AK IV" />
                <AGEGROUP agegroupid="22" agemax="-1" agemin="66" name="offen - Masters AK V" />
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="18" number="18" gender="F" round="TIM">
              <SWIMSTYLE stroke="IMMERSION" technique="DIVE" relaycount="1" distance="100" />
              <FEE value="600" currency="EUR" />
              <HEATS>
                <HEAT heatid="18001" number="1" />
                <HEAT heatid="18002" number="2" />
                <HEAT heatid="18003" number="3" />
                <HEAT heatid="18004" number="4" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="3" agemax="13" agemin="12" name="Sachsen - Altersklasse D">
                  <RANKINGS>
                    <RANKING place="1" resultid="283" />
                    <RANKING place="2" resultid="419" />
                    <RANKING place="3" resultid="493" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="15" agemin="14" name="Sachsen - Altersklasse C">
                  <RANKINGS>
                    <RANKING place="2" resultid="336" />
                    <RANKING place="1" resultid="473" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="17" agemin="16" name="Sachsen - Altersklasse B">
                  <RANKINGS>
                    <RANKING place="2" resultid="299" />
                    <RANKING place="1" resultid="466" />
                    <RANKING place="3" resultid="613" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6" agemax="34" agemin="18" name="Sachsen - Altersklasse A">
                  <RANKINGS>
                    <RANKING place="3" resultid="629" />
                    <RANKING place="2" resultid="636" />
                    <RANKING place="1" resultid="642" />
                    <RANKING place="4" resultid="655" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9" agemax="13" agemin="12" name="offen - Altersklasse D">
                  <RANKINGS>
                    <RANKING place="1" resultid="7" />
                    <RANKING place="5" resultid="131" />
                    <RANKING place="2" resultid="283" />
                    <RANKING place="3" resultid="419" />
                    <RANKING place="4" resultid="493" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10" agemax="15" agemin="14" name="offen - Altersklasse C">
                  <RANKINGS>
                    <RANKING place="4" resultid="33" />
                    <RANKING place="2" resultid="336" />
                    <RANKING place="1" resultid="473" />
                    <RANKING place="3" resultid="667" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11" agemax="17" agemin="16" name="offen - Altersklasse B">
                  <RANKINGS>
                    <RANKING place="2" resultid="16" />
                    <RANKING place="1" resultid="68" />
                    <RANKING place="3" resultid="89" />
                    <RANKING place="7" resultid="299" />
                    <RANKING place="6" resultid="466" />
                    <RANKING place="4" resultid="551" />
                    <RANKING place="8" resultid="613" />
                    <RANKING place="5" resultid="688" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="12" agemax="34" agemin="18" name="offen - Altersklasse A">
                  <RANKINGS>
                    <RANKING place="4" resultid="10" />
                    <RANKING place="3" resultid="72" />
                    <RANKING place="7" resultid="389" />
                    <RANKING place="5" resultid="629" />
                    <RANKING place="2" resultid="636" />
                    <RANKING place="1" resultid="642" />
                    <RANKING place="6" resultid="655" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="13" agemax="44" agemin="35" name="Sachsen - Masters AK I">
                  <RANKINGS>
                    <RANKING place="1" resultid="607" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="14" agemax="45" agemin="36" name="Sachsen - Masters AK II">
                  <RANKINGS>
                    <RANKING place="1" resultid="607" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15" agemax="55" agemin="46" name="Sachsen - Masters AK III" />
                <AGEGROUP agegroupid="16" agemax="65" agemin="56" name="Sachsen - Masters AK IV">
                  <RANKINGS>
                    <RANKING place="1" resultid="359" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="17" agemax="-1" agemin="66" name="Sachsen - Masters AK V" />
                <AGEGROUP agegroupid="18" agemax="44" agemin="35" name="offen - Masters AK I">
                  <RANKINGS>
                    <RANKING place="1" resultid="607" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="19" agemax="45" agemin="36" name="offen - Masters AK II">
                  <RANKINGS>
                    <RANKING place="1" resultid="607" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="20" agemax="55" agemin="46" name="offen - Masters AK III" />
                <AGEGROUP agegroupid="21" agemax="65" agemin="56" name="offen - Masters AK IV">
                  <RANKINGS>
                    <RANKING place="1" resultid="359" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="22" agemax="-1" agemin="66" name="offen - Masters AK V" />
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="19" number="19" gender="M" round="TIM">
              <SWIMSTYLE stroke="IMMERSION" technique="DIVE" relaycount="1" distance="100" />
              <FEE value="600" currency="EUR" />
              <HEATS>
                <HEAT heatid="19001" number="1" />
                <HEAT heatid="19002" number="2" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="3" agemax="13" agemin="12" name="Sachsen - Altersklasse D">
                  <RANKINGS>
                    <RANKING place="1" resultid="424" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="15" agemin="14" name="Sachsen - Altersklasse C" />
                <AGEGROUP agegroupid="5" agemax="17" agemin="16" name="Sachsen - Altersklasse B" />
                <AGEGROUP agegroupid="6" agemax="34" agemin="18" name="Sachsen - Altersklasse A">
                  <RANKINGS>
                    <RANKING place="1" resultid="51" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9" agemax="13" agemin="12" name="offen - Altersklasse D">
                  <RANKINGS>
                    <RANKING place="2" resultid="424" />
                    <RANKING place="1" resultid="718" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10" agemax="15" agemin="14" name="offen - Altersklasse C">
                  <RANKINGS>
                    <RANKING place="1" resultid="25" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11" agemax="17" agemin="16" name="offen - Altersklasse B">
                  <RANKINGS>
                    <RANKING place="1" resultid="218" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="12" agemax="34" agemin="18" name="offen - Altersklasse A">
                  <RANKINGS>
                    <RANKING place="3" resultid="37" />
                    <RANKING place="4" resultid="51" />
                    <RANKING place="1" resultid="138" />
                    <RANKING place="2" resultid="541" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="13" agemax="44" agemin="35" name="Sachsen - Masters AK I" />
                <AGEGROUP agegroupid="14" agemax="45" agemin="36" name="Sachsen - Masters AK II">
                  <RANKINGS>
                    <RANKING place="1" resultid="601" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15" agemax="55" agemin="46" name="Sachsen - Masters AK III">
                  <RANKINGS>
                    <RANKING place="2" resultid="46" />
                    <RANKING place="1" resultid="374" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="16" agemax="65" agemin="56" name="Sachsen - Masters AK IV">
                  <RANKINGS>
                    <RANKING place="1" resultid="57" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="17" agemax="-1" agemin="66" name="Sachsen - Masters AK V">
                  <RANKINGS>
                    <RANKING place="1" resultid="328" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="18" agemax="44" agemin="35" name="offen - Masters AK I" />
                <AGEGROUP agegroupid="19" agemax="45" agemin="36" name="offen - Masters AK II">
                  <RANKINGS>
                    <RANKING place="1" resultid="601" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="20" agemax="55" agemin="46" name="offen - Masters AK III">
                  <RANKINGS>
                    <RANKING place="2" resultid="46" />
                    <RANKING place="1" resultid="374" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="21" agemax="65" agemin="56" name="offen - Masters AK IV">
                  <RANKINGS>
                    <RANKING place="1" resultid="57" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="22" agemax="-1" agemin="66" name="offen - Masters AK V">
                  <RANKINGS>
                    <RANKING place="1" resultid="328" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="20" number="20" gender="F" round="TIM">
              <SWIMSTYLE stroke="SURFACE" relaycount="1" distance="200" />
              <FEE value="600" currency="EUR" />
              <HEATS>
                <HEAT heatid="20001" number="1" />
                <HEAT heatid="20002" number="2" />
                <HEAT heatid="20003" number="3" />
                <HEAT heatid="20004" number="4" />
                <HEAT heatid="20005" number="5" />
                <HEAT heatid="20006" number="6" />
                <HEAT heatid="20007" number="7" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="10" agemin="7" name="Sachsen - Altersklasse F">
                  <RANKINGS>
                    <RANKING place="2" resultid="469" />
                    <RANKING place="1" resultid="502" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2" agemax="11" agemin="11" name="Sachsen - Altersklasse E">
                  <RANKINGS>
                    <RANKING place="1" resultid="350" />
                    <RANKING place="2" resultid="381" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3" agemax="13" agemin="12" name="Sachsen - Altersklasse D">
                  <RANKINGS>
                    <RANKING place="4" resultid="290" />
                    <RANKING place="5" resultid="378" />
                    <RANKING place="3" resultid="396" />
                    <RANKING place="1" resultid="400" />
                    <RANKING place="2" resultid="420" />
                    <RANKING place="6" resultid="457" />
                    <RANKING place="7" resultid="480" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="15" agemin="14" name="Sachsen - Altersklasse C">
                  <RANKINGS>
                    <RANKING place="2" resultid="296" />
                    <RANKING place="4" resultid="371" />
                    <RANKING place="3" resultid="460" />
                    <RANKING place="1" resultid="708" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="17" agemin="16" name="Sachsen - Altersklasse B">
                  <RANKINGS>
                    <RANKING place="2" resultid="63" />
                    <RANKING place="3" resultid="591" />
                    <RANKING place="1" resultid="621" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6" agemax="34" agemin="18" name="Sachsen - Altersklasse A">
                  <RANKINGS>
                    <RANKING place="4" resultid="415" />
                    <RANKING place="3" resultid="445" />
                    <RANKING place="1" resultid="637" />
                    <RANKING place="2" resultid="656" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7" agemax="10" agemin="7" name="offen - Altersklasse F">
                  <RANKINGS>
                    <RANKING place="4" resultid="99" />
                    <RANKING place="1" resultid="103" />
                    <RANKING place="3" resultid="469" />
                    <RANKING place="2" resultid="502" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8" agemax="11" agemin="11" name="offen - Altersklasse E">
                  <RANKINGS>
                    <RANKING place="1" resultid="350" />
                    <RANKING place="2" resultid="381" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9" agemax="13" agemin="12" name="offen - Altersklasse D">
                  <RANKINGS>
                    <RANKING place="9" resultid="96" />
                    <RANKING place="6" resultid="290" />
                    <RANKING place="7" resultid="378" />
                    <RANKING place="5" resultid="396" />
                    <RANKING place="2" resultid="400" />
                    <RANKING place="3" resultid="420" />
                    <RANKING place="8" resultid="457" />
                    <RANKING place="10" resultid="480" />
                    <RANKING place="1" resultid="663" />
                    <RANKING place="4" resultid="672" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10" agemax="15" agemin="14" name="offen - Altersklasse C">
                  <RANKINGS>
                    <RANKING place="7" resultid="34" />
                    <RANKING place="3" resultid="296" />
                    <RANKING place="8" resultid="371" />
                    <RANKING place="4" resultid="460" />
                    <RANKING place="1" resultid="560" />
                    <RANKING place="5" resultid="668" />
                    <RANKING place="6" resultid="696" />
                    <RANKING place="2" resultid="708" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11" agemax="17" agemin="16" name="offen - Altersklasse B">
                  <RANKINGS>
                    <RANKING place="6" resultid="63" />
                    <RANKING place="1" resultid="148" />
                    <RANKING place="3" resultid="243" />
                    <RANKING place="4" resultid="254" />
                    <RANKING place="2" resultid="566" />
                    <RANKING place="7" resultid="591" />
                    <RANKING place="5" resultid="621" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="12" agemax="34" agemin="18" name="offen - Altersklasse A">
                  <RANKINGS>
                    <RANKING place="2" resultid="73" />
                    <RANKING place="5" resultid="113" />
                    <RANKING place="7" resultid="415" />
                    <RANKING place="6" resultid="445" />
                    <RANKING place="1" resultid="546" />
                    <RANKING place="3" resultid="637" />
                    <RANKING place="4" resultid="656" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="13" agemax="44" agemin="35" name="Sachsen - Masters AK I" />
                <AGEGROUP agegroupid="14" agemax="45" agemin="36" name="Sachsen - Masters AK II" />
                <AGEGROUP agegroupid="15" agemax="55" agemin="46" name="Sachsen - Masters AK III" />
                <AGEGROUP agegroupid="16" agemax="65" agemin="56" name="Sachsen - Masters AK IV" />
                <AGEGROUP agegroupid="17" agemax="-1" agemin="66" name="Sachsen - Masters AK V" />
                <AGEGROUP agegroupid="18" agemax="44" agemin="35" name="offen - Masters AK I" />
                <AGEGROUP agegroupid="19" agemax="45" agemin="36" name="offen - Masters AK II" />
                <AGEGROUP agegroupid="20" agemax="55" agemin="46" name="offen - Masters AK III">
                  <RANKINGS>
                    <RANKING place="1" resultid="200" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="21" agemax="65" agemin="56" name="offen - Masters AK IV">
                  <RANKINGS>
                    <RANKING place="1" resultid="704" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="22" agemax="-1" agemin="66" name="offen - Masters AK V" />
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="21" number="21" gender="M" round="TIM">
              <SWIMSTYLE stroke="SURFACE" relaycount="1" distance="200" />
              <FEE value="600" currency="EUR" />
              <HEATS>
                <HEAT heatid="21001" number="1" />
                <HEAT heatid="21002" number="2" />
                <HEAT heatid="21003" number="3" />
                <HEAT heatid="21004" number="4" />
                <HEAT heatid="21005" number="5" />
                <HEAT heatid="21006" number="6" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="10" agemin="7" name="Sachsen - Altersklasse F">
                  <RANKINGS>
                    <RANKING place="2" resultid="275" />
                    <RANKING place="4" resultid="286" />
                    <RANKING place="5" resultid="332" />
                    <RANKING place="3" resultid="353" />
                    <RANKING place="1" resultid="356" />
                    <RANKING place="6" resultid="384" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2" agemax="11" agemin="11" name="Sachsen - Altersklasse E">
                  <RANKINGS>
                    <RANKING place="1" resultid="486" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3" agemax="13" agemin="12" name="Sachsen - Altersklasse D">
                  <RANKINGS>
                    <RANKING place="1" resultid="425" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="15" agemin="14" name="Sachsen - Altersklasse C">
                  <RANKINGS>
                    <RANKING place="2" resultid="279" />
                    <RANKING place="3" resultid="306" />
                    <RANKING place="1" resultid="320" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="17" agemin="16" name="Sachsen - Altersklasse B">
                  <RANKINGS>
                    <RANKING place="2" resultid="412" />
                    <RANKING place="1" resultid="440" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6" agemax="34" agemin="18" name="Sachsen - Altersklasse A" />
                <AGEGROUP agegroupid="7" agemax="10" agemin="7" name="offen - Altersklasse F">
                  <RANKINGS>
                    <RANKING place="1" resultid="127" />
                    <RANKING place="9" resultid="134" />
                    <RANKING place="2" resultid="142" />
                    <RANKING place="4" resultid="275" />
                    <RANKING place="6" resultid="286" />
                    <RANKING place="7" resultid="332" />
                    <RANKING place="5" resultid="353" />
                    <RANKING place="3" resultid="356" />
                    <RANKING place="8" resultid="384" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8" agemax="11" agemin="11" name="offen - Altersklasse E">
                  <RANKINGS>
                    <RANKING place="2" resultid="146" />
                    <RANKING place="3" resultid="265" />
                    <RANKING place="1" resultid="486" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9" agemax="13" agemin="12" name="offen - Altersklasse D">
                  <RANKINGS>
                    <RANKING place="7" resultid="221" />
                    <RANKING place="2" resultid="232" />
                    <RANKING place="5" resultid="236" />
                    <RANKING place="6" resultid="262" />
                    <RANKING place="4" resultid="425" />
                    <RANKING place="8" resultid="680" />
                    <RANKING place="3" resultid="684" />
                    <RANKING place="1" resultid="719" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10" agemax="15" agemin="14" name="offen - Altersklasse C">
                  <RANKINGS>
                    <RANKING place="3" resultid="22" />
                    <RANKING place="1" resultid="26" />
                    <RANKING place="4" resultid="258" />
                    <RANKING place="7" resultid="279" />
                    <RANKING place="8" resultid="306" />
                    <RANKING place="2" resultid="320" />
                    <RANKING place="5" resultid="676" />
                    <RANKING place="6" resultid="714" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11" agemax="17" agemin="16" name="offen - Altersklasse B">
                  <RANKINGS>
                    <RANKING place="3" resultid="412" />
                    <RANKING place="2" resultid="440" />
                    <RANKING place="4" resultid="538" />
                    <RANKING place="5" resultid="574" />
                    <RANKING place="1" resultid="692" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="12" agemax="34" agemin="18" name="offen - Altersklasse A">
                  <RANKINGS>
                    <RANKING place="1" resultid="570" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="13" agemax="44" agemin="35" name="Sachsen - Masters AK I">
                  <RANKINGS>
                    <RANKING place="1" resultid="587" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="14" agemax="45" agemin="36" name="Sachsen - Masters AK II">
                  <RANKINGS>
                    <RANKING place="1" resultid="587" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15" agemax="55" agemin="46" name="Sachsen - Masters AK III">
                  <RANKINGS>
                    <RANKING place="2" resultid="47" />
                    <RANKING place="1" resultid="520" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="16" agemax="65" agemin="56" name="Sachsen - Masters AK IV">
                  <RANKINGS>
                    <RANKING place="2" resultid="58" />
                    <RANKING place="3" resultid="368" />
                    <RANKING place="1" resultid="531" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="17" agemax="-1" agemin="66" name="Sachsen - Masters AK V" />
                <AGEGROUP agegroupid="18" agemax="44" agemin="35" name="offen - Masters AK I">
                  <RANKINGS>
                    <RANKING place="1" resultid="587" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="19" agemax="45" agemin="36" name="offen - Masters AK II">
                  <RANKINGS>
                    <RANKING place="1" resultid="587" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="20" agemax="55" agemin="46" name="offen - Masters AK III">
                  <RANKINGS>
                    <RANKING place="2" resultid="47" />
                    <RANKING place="3" resultid="119" />
                    <RANKING place="1" resultid="520" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="21" agemax="65" agemin="56" name="offen - Masters AK IV">
                  <RANKINGS>
                    <RANKING place="2" resultid="58" />
                    <RANKING place="3" resultid="368" />
                    <RANKING place="1" resultid="531" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="22" agemax="-1" agemin="66" name="offen - Masters AK V" />
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="22" number="22" gender="F" round="TIM">
              <SWIMSTYLE stroke="IMMERSION" technique="DIVE" relaycount="1" distance="400" />
              <FEE value="600" currency="EUR" />
              <HEATS>
                <HEAT heatid="22001" number="1" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="3" agemax="13" agemin="12" name="Sachsen - Altersklasse D" />
                <AGEGROUP agegroupid="4" agemax="15" agemin="14" name="Sachsen - Altersklasse C">
                  <RANKINGS>
                    <RANKING place="1" resultid="705" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="17" agemin="16" name="Sachsen - Altersklasse B" />
                <AGEGROUP agegroupid="6" agemax="34" agemin="18" name="Sachsen - Altersklasse A">
                  <RANKINGS>
                    <RANKING place="2" resultid="650" />
                    <RANKING place="1" resultid="657" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9" agemax="13" agemin="12" name="offen - Altersklasse D" />
                <AGEGROUP agegroupid="10" agemax="15" agemin="14" name="offen - Altersklasse C">
                  <RANKINGS>
                    <RANKING place="1" resultid="705" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11" agemax="17" agemin="16" name="offen - Altersklasse B">
                  <RANKINGS>
                    <RANKING place="1" resultid="17" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="12" agemax="34" agemin="18" name="offen - Altersklasse A">
                  <RANKINGS>
                    <RANKING place="1" resultid="11" />
                    <RANKING place="3" resultid="30" />
                    <RANKING place="4" resultid="650" />
                    <RANKING place="2" resultid="657" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="13" agemax="44" agemin="35" name="Sachsen - Masters AK I" />
                <AGEGROUP agegroupid="14" agemax="45" agemin="36" name="Sachsen - Masters AK II" />
                <AGEGROUP agegroupid="15" agemax="55" agemin="46" name="Sachsen - Masters AK III" />
                <AGEGROUP agegroupid="16" agemax="65" agemin="56" name="Sachsen - Masters AK IV">
                  <RANKINGS>
                    <RANKING place="1" resultid="360" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="17" agemax="-1" agemin="66" name="Sachsen - Masters AK V" />
                <AGEGROUP agegroupid="18" agemax="44" agemin="35" name="offen - Masters AK I" />
                <AGEGROUP agegroupid="19" agemax="45" agemin="36" name="offen - Masters AK II" />
                <AGEGROUP agegroupid="20" agemax="55" agemin="46" name="offen - Masters AK III" />
                <AGEGROUP agegroupid="21" agemax="65" agemin="56" name="offen - Masters AK IV">
                  <RANKINGS>
                    <RANKING place="1" resultid="360" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="22" agemax="-1" agemin="66" name="offen - Masters AK V" />
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="23" number="23" gender="M" round="TIM">
              <SWIMSTYLE stroke="IMMERSION" technique="DIVE" relaycount="1" distance="400" />
              <FEE value="600" currency="EUR" />
              <HEATS>
                <HEAT heatid="23001" number="1" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="3" agemax="13" agemin="12" name="Sachsen - Altersklasse D" />
                <AGEGROUP agegroupid="4" agemax="15" agemin="14" name="Sachsen - Altersklasse C" />
                <AGEGROUP agegroupid="5" agemax="17" agemin="16" name="Sachsen - Altersklasse B" />
                <AGEGROUP agegroupid="6" agemax="34" agemin="18" name="Sachsen - Altersklasse A">
                  <RANKINGS>
                    <RANKING place="1" resultid="302" />
                    <RANKING place="2" resultid="624" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9" agemax="13" agemin="12" name="offen - Altersklasse D" />
                <AGEGROUP agegroupid="10" agemax="15" agemin="14" name="offen - Altersklasse C" />
                <AGEGROUP agegroupid="11" agemax="17" agemin="16" name="offen - Altersklasse B">
                  <RANKINGS>
                    <RANKING place="1" resultid="575" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="12" agemax="34" agemin="18" name="offen - Altersklasse A">
                  <RANKINGS>
                    <RANKING place="1" resultid="3" />
                    <RANKING place="3" resultid="38" />
                    <RANKING place="2" resultid="302" />
                    <RANKING place="4" resultid="624" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="13" agemax="44" agemin="35" name="Sachsen - Masters AK I" />
                <AGEGROUP agegroupid="14" agemax="45" agemin="36" name="Sachsen - Masters AK II" />
                <AGEGROUP agegroupid="15" agemax="55" agemin="46" name="Sachsen - Masters AK III" />
                <AGEGROUP agegroupid="16" agemax="65" agemin="56" name="Sachsen - Masters AK IV">
                  <RANKINGS>
                    <RANKING place="1" resultid="59" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="17" agemax="-1" agemin="66" name="Sachsen - Masters AK V" />
                <AGEGROUP agegroupid="18" agemax="44" agemin="35" name="offen - Masters AK I" />
                <AGEGROUP agegroupid="19" agemax="45" agemin="36" name="offen - Masters AK II" />
                <AGEGROUP agegroupid="20" agemax="55" agemin="46" name="offen - Masters AK III" />
                <AGEGROUP agegroupid="21" agemax="65" agemin="56" name="offen - Masters AK IV">
                  <RANKINGS>
                    <RANKING place="1" resultid="59" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="22" agemax="-1" agemin="66" name="offen - Masters AK V" />
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="24" number="24" gender="F" round="TIM">
              <SWIMSTYLE stroke="SURFACE" relaycount="4" distance="100" />
              <FEE value="800" currency="EUR" />
              <HEATS>
                <HEAT heatid="24001" number="1" />
                <HEAT heatid="24002" number="2" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="14" agemin="7" name="Sachsen - Kategorie A">
                  <RANKINGS>
                    <RANKING place="1" resultid="322" />
                    <RANKING place="2" resultid="431" />
                    <RANKING place="3" resultid="647" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2" agemax="18" agemin="15" name="Sachsen - Kategorie B">
                  <RANKINGS>
                    <RANKING place="1" resultid="270" />
                    <RANKING place="2" resultid="646" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3" agemax="-1" agemin="19" name="Sachsen - Kategorie A">
                  <RANKINGS>
                    <RANKING place="1" resultid="427" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="14" agemin="7" name="offen - Kategorie A">
                  <RANKINGS>
                    <RANKING place="2" resultid="322" />
                    <RANKING place="3" resultid="431" />
                    <RANKING place="4" resultid="647" />
                    <RANKING place="1" resultid="659" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="18" agemin="15" name="offen - Kategorie B">
                  <RANKINGS>
                    <RANKING place="2" resultid="270" />
                    <RANKING place="1" resultid="534" />
                    <RANKING place="3" resultid="646" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6" agemax="-1" agemin="19" name="offen - Kategorie A">
                  <RANKINGS>
                    <RANKING place="1" resultid="427" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7" agemax="-1" agemin="176" easy.ak="176" calculate="TOTAL" name="Sachsen - Masters A" />
                <AGEGROUP agegroupid="8" agemax="-1" agemin="399" easy.ak="399" calculate="TOTAL" name="Sachsen - Masters B" />
                <AGEGROUP agegroupid="9" agemax="-1" agemin="176" easy.ak="176" calculate="TOTAL" name="offen - Masters A" />
                <AGEGROUP agegroupid="10" agemax="-1" agemin="399" easy.ak="399" calculate="TOTAL" name="offen - Masters B" />
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="25" number="25" gender="M" round="TIM">
              <SWIMSTYLE stroke="SURFACE" relaycount="4" distance="100" />
              <FEE value="800" currency="EUR" />
              <HEATS>
                <HEAT heatid="25001" number="1" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="14" agemin="7" name="Sachsen - Kategorie A" />
                <AGEGROUP agegroupid="2" agemax="18" agemin="15" name="Sachsen - Kategorie B">
                  <RANKINGS>
                    <RANKING place="1" resultid="268" />
                    <RANKING place="2" resultid="429" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3" agemax="-1" agemin="19" name="Sachsen - Kategorie A">
                  <RANKINGS>
                    <RANKING place="1" resultid="428" />
                    <RANKING place="3" resultid="503" />
                    <RANKING place="2" resultid="581" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="14" agemin="7" name="offen - Kategorie A" />
                <AGEGROUP agegroupid="5" agemax="18" agemin="15" name="offen - Kategorie B">
                  <RANKINGS>
                    <RANKING place="1" resultid="268" />
                    <RANKING place="2" resultid="429" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6" agemax="-1" agemin="19" name="offen - Kategorie A">
                  <RANKINGS>
                    <RANKING place="1" resultid="428" />
                    <RANKING place="4" resultid="503" />
                    <RANKING place="2" resultid="532" />
                    <RANKING place="3" resultid="581" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7" agemax="-1" agemin="176" easy.ak="176" calculate="TOTAL" name="Sachsen - Masters A">
                  <RANKINGS>
                    <RANKING place="1" resultid="503" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8" agemax="-1" agemin="399" easy.ak="399" calculate="TOTAL" name="Sachsen - Masters B" />
                <AGEGROUP agegroupid="9" agemax="-1" agemin="176" easy.ak="176" calculate="TOTAL" name="offen - Masters A">
                  <RANKINGS>
                    <RANKING place="1" resultid="503" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10" agemax="-1" agemin="399" easy.ak="399" calculate="TOTAL" name="offen - Masters B" />
              </AGEGROUPS>
            </EVENT>
          </EVENTS>
        </SESSION>
      </SESSIONS>
      <CLUBS>
        <CLUB name="1. Chemnitzer Tauchverein e.V." nation="GER" region="20" code="0">
          <ATHLETES>
            <ATHLETE athleteid="104" birthdate="2013-01-01" gender="M" lastname="Münzner" firstname="Alfred" license="0">
              <RESULTS>
                <RESULT resultid="273" eventid="2" swimtime="00:06:12.90" reactiontime="+80" lane="7" heatid="2002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:23.39" />
                    <SPLIT distance="200" swimtime="00:02:59.63" />
                    <SPLIT distance="300" swimtime="00:04:38.48" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="274" eventid="15" swimtime="00:00:33.36" lane="2" heatid="15004" />
                <RESULT resultid="275" eventid="21" swimtime="00:03:00.98" reactiontime="+93" lane="2" heatid="21002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:25.71" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="105" birthdate="2009-01-01" gender="M" lastname="Müller" firstname="Alwin" license="0">
              <RESULTS>
                <RESULT resultid="276" eventid="6" swimtime="00:00:27.60" lane="5" heatid="6001" />
                <RESULT resultid="277" eventid="8" swimtime="00:01:05.54" reactiontime="+84" lane="4" heatid="8004" />
                <RESULT resultid="278" eventid="15" swimtime="00:00:28.66" lane="6" heatid="15005" />
                <RESULT resultid="279" eventid="21" swimtime="00:02:26.64" reactiontime="+87" lane="8" heatid="21004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:10.00" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="106" birthdate="2010-01-01" gender="F" lastname="Schwarzer" firstname="Angelina Sophie" license="0">
              <RESULTS>
                <RESULT resultid="280" eventid="1" swimtime="00:04:38.71" reactiontime="+96" lane="8" heatid="1003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:59.83" />
                    <SPLIT distance="200" swimtime="00:02:13.21" />
                    <SPLIT distance="300" swimtime="00:03:28.71" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="281" eventid="7" swimtime="00:00:58.33" lane="7" heatid="7007" />
                <RESULT resultid="282" eventid="14" swimtime="00:00:26.30" lane="3" heatid="14007" />
                <RESULT resultid="283" eventid="18" swimtime="00:01:00.79" lane="7" heatid="18002" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="107" birthdate="2013-01-01" gender="M" lastname="Schiller" firstname="Ben" license="0">
              <RESULTS>
                <RESULT resultid="284" eventid="8" swimtime="00:01:23.36" reactiontime="+95" lane="6" heatid="8002" />
                <RESULT resultid="285" eventid="15" swimtime="00:00:37.49" lane="2" heatid="15002" />
                <RESULT resultid="286" eventid="21" swimtime="00:03:13.43" reactiontime="+99" lane="8" heatid="21002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:30.45" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="108" birthdate="2010-01-01" gender="F" lastname="Siegert" firstname="Emilia" license="0">
              <RESULTS>
                <RESULT resultid="287" eventid="3" swimtime="00:00:31.50" lane="3" heatid="3001" />
                <RESULT resultid="288" eventid="7" swimtime="00:01:04.05" reactiontime="+97" lane="8" heatid="7006" />
                <RESULT resultid="289" eventid="14" swimtime="00:00:30.47" lane="1" heatid="14007" />
                <RESULT resultid="290" eventid="20" swimtime="00:02:24.31" reactiontime="+93" lane="5" heatid="20004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:11.20" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="109" birthdate="2011-01-01" gender="F" lastname="Nisch" firstname="Hanna Maria" license="0">
              <RESULTS>
                <RESULT resultid="291" eventid="1" swimtime="00:04:47.59" reactiontime="+97" lane="1" heatid="1003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:08.31" />
                    <SPLIT distance="200" swimtime="00:02:23.16" />
                    <SPLIT distance="300" swimtime="00:03:39.06" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="292" eventid="7" swimtime="00:01:01.70" lane="2" heatid="7006" />
                <RESULT resultid="293" eventid="18" status="DSQ" swimtime="00:00:00.00" lane="2" heatid="18002" comment="Gesicht aus dem Wasser bei 40 Meter." />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="110" birthdate="2008-01-01" gender="F" lastname="Franke" firstname="Jenny" license="0">
              <RESULTS>
                <RESULT resultid="294" eventid="5" swimtime="00:00:21.71" lane="8" heatid="5003" />
                <RESULT resultid="295" eventid="14" swimtime="00:00:22.84" lane="5" heatid="14008" />
                <RESULT resultid="296" eventid="20" swimtime="00:01:57.64" reactiontime="+98" lane="5" heatid="20005">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:56.52" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="111" birthdate="2007-01-01" gender="F" lastname="Ullrich" firstname="Johanna Hermine" license="0">
              <RESULTS>
                <RESULT resultid="297" eventid="5" swimtime="00:00:24.08" lane="2" heatid="5002" />
                <RESULT resultid="298" eventid="9" swimtime="00:08:55.21" reactiontime="+81" lane="1" heatid="9002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:00.27" />
                    <SPLIT distance="200" swimtime="00:02:08.08" />
                    <SPLIT distance="300" swimtime="00:03:15.80" />
                    <SPLIT distance="400" swimtime="00:04:24.82" />
                    <SPLIT distance="500" swimtime="00:05:33.59" />
                    <SPLIT distance="600" swimtime="00:06:42.81" />
                    <SPLIT distance="700" swimtime="00:07:52.74" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="299" eventid="18" swimtime="00:00:57.37" lane="8" heatid="18003" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="112" birthdate="2005-01-01" gender="M" lastname="Porges" firstname="Marcel" license="0">
              <RESULTS>
                <RESULT resultid="300" eventid="6" swimtime="00:00:16.25" lane="5" heatid="6004" />
                <RESULT resultid="301" eventid="15" swimtime="00:00:17.69" lane="6" heatid="15009" />
                <RESULT resultid="302" eventid="23" swimtime="00:03:18.73" lane="5" heatid="23001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:45.81" />
                    <SPLIT distance="200" swimtime="00:01:36.39" />
                    <SPLIT distance="300" swimtime="00:02:28.27" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="113" birthdate="2009-01-01" gender="M" lastname="Elle" firstname="Simon" license="0">
              <RESULTS>
                <RESULT resultid="303" eventid="4" swimtime="00:00:37.64" lane="6" heatid="4001" />
                <RESULT resultid="304" eventid="8" swimtime="00:01:15.99" reactiontime="+72" lane="2" heatid="8003" />
                <RESULT resultid="305" eventid="15" swimtime="00:00:33.71" lane="8" heatid="15004" />
                <RESULT resultid="306" eventid="21" swimtime="00:02:37.56" reactiontime="+82" lane="3" heatid="21002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:13.48" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="114" birthdate="2013-01-01" gender="F" lastname="Wende" firstname="Sophia" license="0">
              <RESULTS>
                <RESULT resultid="307" eventid="1" status="DNS" swimtime="00:00:00.00" lane="5" heatid="1001" />
                <RESULT resultid="308" eventid="14" status="DNS" swimtime="00:00:00.00" lane="4" heatid="14002" />
                <RESULT resultid="309" eventid="20" status="DNS" swimtime="00:00:00.00" lane="2" heatid="20002" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="115" birthdate="2010-01-01" gender="F" lastname="Bluhm" firstname="Suna" license="0">
              <RESULTS>
                <RESULT resultid="310" eventid="3" status="DNS" swimtime="00:00:00.00" lane="7" heatid="3001" />
                <RESULT resultid="311" eventid="7" status="DNS" swimtime="00:00:00.00" lane="7" heatid="7005" />
                <RESULT resultid="312" eventid="14" status="DNS" swimtime="00:00:00.00" lane="2" heatid="14005" />
                <RESULT resultid="313" eventid="20" status="DNS" swimtime="00:00:00.00" lane="8" heatid="20004" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="116" birthdate="2012-01-01" gender="M" lastname="Ilianyi" firstname="Yan" license="0">
              <RESULTS>
                <RESULT resultid="314" eventid="8" swimtime="00:01:25.18" reactiontime="+65" lane="3" heatid="8002" />
                <RESULT resultid="315" eventid="15" swimtime="00:00:39.32" lane="1" heatid="15003" />
                <RESULT resultid="316" eventid="21" status="DSQ" swimtime="00:03:39.18" lane="1" heatid="21002" comment="Aufgegeben nach 80 Meter.">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:52.42" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="117" birthdate="2009-01-01" gender="M" lastname="Hans" firstname="Yannick" license="0">
              <RESULTS>
                <RESULT resultid="317" eventid="6" swimtime="00:00:23.23" lane="6" heatid="6002" />
                <RESULT resultid="318" eventid="8" swimtime="00:00:54.59" reactiontime="+95" lane="5" heatid="8006" />
                <RESULT resultid="319" eventid="15" swimtime="00:00:24.84" lane="8" heatid="15007" />
                <RESULT resultid="320" eventid="21" swimtime="00:01:59.82" reactiontime="+96" lane="2" heatid="21005">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:58.88" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY number="1" gender="M" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="268" eventid="25" swimtime="00:04:05.92" lane="2" heatid="25001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:41.20" />
                    <SPLIT distance="200" swimtime="00:01:46.98" />
                    <SPLIT distance="300" swimtime="00:03:11.45" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="112" number="1" />
                    <RELAYPOSITION athleteid="105" number="2" />
                    <RELAYPOSITION athleteid="104" number="3" />
                    <RELAYPOSITION athleteid="117" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="2" gender="X" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="269" eventid="13" swimtime="00:01:29.70" lane="6" heatid="13002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:47.02" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="117" number="1" />
                    <RELAYPOSITION athleteid="110" number="2" />
                    <RELAYPOSITION athleteid="111" number="3" />
                    <RELAYPOSITION athleteid="112" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="3" gender="F" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="270" eventid="24" swimtime="00:03:49.64" lane="6" heatid="24002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:01.09" />
                    <SPLIT distance="200" swimtime="00:01:57.71" />
                    <SPLIT distance="300" swimtime="00:02:58.74" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="109" number="1" />
                    <RELAYPOSITION athleteid="111" number="2" />
                    <RELAYPOSITION athleteid="106" number="3" />
                    <RELAYPOSITION athleteid="110" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="4" gender="X" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="271" eventid="13" status="DSQ" swimtime="00:02:00.15" lane="8" heatid="13002" comment="4. Starter: Falsche Ausrüstung.">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:56.33" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="108" number="1" />
                    <RELAYPOSITION athleteid="109" number="2" />
                    <RELAYPOSITION athleteid="105" number="3" />
                    <RELAYPOSITION athleteid="104" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="5" gender="X" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="272" eventid="13" swimtime="00:02:17.50" lane="6" heatid="13001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:13.08" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="113" number="1" />
                    <RELAYPOSITION athleteid="107" number="2" />
                    <RELAYPOSITION athleteid="116" number="3" />
                    <RELAYPOSITION athleteid="106" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB name="Berliner TSC e.V." nation="GER" region="21" code="304088">
          <ATHLETES>
            <ATHLETE athleteid="50" birthdate="2007-01-01" gender="F" lastname="Manthey" firstname="Maxime" license="123">
              <RESULTS>
                <RESULT resultid="147" eventid="14" swimtime="00:00:20.43" lane="7" heatid="14011" />
                <RESULT resultid="148" eventid="20" swimtime="00:01:41.84" reactiontime="+84" lane="2" heatid="20007">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:47.94" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="DJK VfR Mülheim Saarn" nation="GER" region="28" code="8006000">
          <ATHLETES>
            <ATHLETE athleteid="1" birthdate="2005-01-01" gender="M" lastname="Bieler" firstname="Phil Jason" license="0">
              <RESULTS>
                <RESULT resultid="1" eventid="10" swimtime="00:07:05.86" reactiontime="+97" lane="5" heatid="10001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:47.59" />
                    <SPLIT distance="200" swimtime="00:01:40.81" />
                    <SPLIT distance="300" swimtime="00:02:34.98" />
                    <SPLIT distance="400" swimtime="00:03:29.37" />
                    <SPLIT distance="500" swimtime="00:04:24.66" />
                    <SPLIT distance="600" swimtime="00:05:20.30" />
                    <SPLIT distance="700" swimtime="00:06:14.00" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="2" eventid="17" swimtime="00:13:49.10" reactiontime="+98" lane="4" heatid="17001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:48.30" />
                    <SPLIT distance="200" swimtime="00:01:43.16" />
                    <SPLIT distance="300" swimtime="00:02:39.30" />
                    <SPLIT distance="400" swimtime="00:03:35.19" />
                    <SPLIT distance="500" swimtime="00:04:31.31" />
                    <SPLIT distance="600" swimtime="00:05:27.54" />
                    <SPLIT distance="700" swimtime="00:06:23.46" />
                    <SPLIT distance="800" swimtime="00:07:20.75" />
                    <SPLIT distance="900" swimtime="00:08:16.86" />
                    <SPLIT distance="1000" swimtime="00:09:12.08" />
                    <SPLIT distance="1100" swimtime="00:10:08.65" />
                    <SPLIT distance="1200" swimtime="00:11:05.66" />
                    <SPLIT distance="1300" swimtime="00:12:02.91" />
                    <SPLIT distance="1400" swimtime="00:12:58.24" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="3" eventid="23" swimtime="00:03:12.39" lane="4" heatid="23001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:44.48" />
                    <SPLIT distance="200" swimtime="00:01:33.89" />
                    <SPLIT distance="300" swimtime="00:02:24.28" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="2" birthdate="2010-01-01" gender="F" lastname="Lazarenko" firstname="Valeria" license="0">
              <RESULTS>
                <RESULT resultid="4" eventid="3" swimtime="00:00:21.81" lane="5" heatid="3001" />
                <RESULT resultid="5" eventid="9" swimtime="00:08:54.48" reactiontime="+98" lane="7" heatid="9002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:01.54" />
                    <SPLIT distance="200" swimtime="00:02:09.45" />
                    <SPLIT distance="300" swimtime="00:03:17.48" />
                    <SPLIT distance="400" swimtime="00:04:27.01" />
                    <SPLIT distance="500" swimtime="00:05:37.08" />
                    <SPLIT distance="600" swimtime="00:06:46.68" />
                    <SPLIT distance="700" swimtime="00:07:53.38" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="6" eventid="14" swimtime="00:00:23.01" lane="1" heatid="14009" />
                <RESULT resultid="7" eventid="18" swimtime="00:00:50.25" lane="3" heatid="18002" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="Landestauchsportverband Sachsen" nation="GER" region="20" code="99">
          <ATHLETES>
            <ATHLETE athleteid="255" birthdate="2011-01-01" gender="M" lastname="Becker." firstname="Pepe" license="0" />
            <ATHLETE athleteid="256" birthdate="2011-01-01" gender="M" lastname="Schönherr." firstname="Nina" license="0" />
            <ATHLETE athleteid="257" birthdate="2011-01-01" gender="M" lastname="Hönisch." firstname="Ida" license="0" />
            <ATHLETE athleteid="258" birthdate="2010-01-01" gender="M" lastname="Berger." firstname="Lene" license="0" />
            <ATHLETE athleteid="259" birthdate="2006-01-01" gender="M" lastname="Loßner." firstname="Niklas" license="0" />
            <ATHLETE athleteid="260" birthdate="2009-01-01" gender="M" lastname="Batiuk." firstname="Mykyta" license="0" />
            <ATHLETE athleteid="261" birthdate="2008-01-01" gender="F" lastname="Kulchyska." firstname="Polina" license="0" />
            <ATHLETE athleteid="262" birthdate="2008-01-01" gender="F" lastname="Horenok." firstname="Polina" license="0" />
            <ATHLETE athleteid="298" birthdate="2006-01-01" gender="M" lastname="Noack." firstname="Christopher" license="0" />
            <ATHLETE athleteid="299" birthdate="1994-01-01" gender="M" lastname="Poschart." firstname="Max" license="0" />
          </ATHLETES>
          <RELAYS>
            <RELAY number="1" gender="F" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="392" eventid="24" status="WDR" swimtime="00:00:00.00" lane="3" heatid="24001" />
              </RESULTS>
            </RELAY>
            <RELAY number="2" gender="M" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="581" eventid="25" swimtime="00:02:55.34" lane="7" heatid="25001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:34.68" />
                    <SPLIT distance="200" swimtime="00:01:29.68" />
                    <SPLIT distance="300" swimtime="00:02:08.49" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="299" number="1" />
                    <RELAYPOSITION athleteid="298" number="2" />
                    <RELAYPOSITION athleteid="259" number="3" />
                    <RELAYPOSITION athleteid="260" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="3" gender="X" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="582" eventid="13" swimtime="00:01:53.11" lane="7" heatid="13001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:55.40" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="255" number="1" />
                    <RELAYPOSITION athleteid="256" number="2" />
                    <RELAYPOSITION athleteid="257" number="3" />
                    <RELAYPOSITION athleteid="258" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB name="SC DHfK Leipzig Flossenschwimmen" nation="GER" region="20" code="0">
          <ATHLETES>
            <ATHLETE athleteid="158" birthdate="2008-01-01" gender="M" lastname="Berger" firstname="Alex Michael" license="0">
              <RESULTS>
                <RESULT resultid="433" eventid="2" swimtime="00:04:00.39" reactiontime="+91" lane="1" heatid="2004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:55.77" />
                    <SPLIT distance="200" swimtime="00:01:59.91" />
                    <SPLIT distance="300" swimtime="00:03:02.80" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="434" eventid="8" swimtime="00:00:47.42" reactiontime="+99" lane="2" heatid="8007" />
                <RESULT resultid="435" eventid="15" status="DNS" swimtime="00:00:00.00" lane="8" heatid="15008" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="159" birthdate="2013-01-01" gender="M" lastname="Beyer" firstname="Arved" license="0">
              <RESULTS>
                <RESULT resultid="709" eventid="8" swimtime="00:01:30.01" lane="2" heatid="8002" />
                <RESULT resultid="436" eventid="15" swimtime="00:00:39.51" lane="6" heatid="15002" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="160" birthdate="2007-01-01" gender="M" lastname="Schoodt" firstname="Ben Joseph" license="2944">
              <RESULTS>
                <RESULT resultid="437" eventid="6" swimtime="00:00:16.86" lane="6" heatid="6004" />
                <RESULT resultid="438" eventid="8" swimtime="00:00:42.97" reactiontime="+94" lane="1" heatid="8008" />
                <RESULT resultid="439" eventid="15" swimtime="00:00:19.30" lane="2" heatid="15009" />
                <RESULT resultid="440" eventid="21" swimtime="00:01:37.28" reactiontime="+93" lane="6" heatid="21006">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:47.22" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="161" birthdate="2014-01-01" gender="F" lastname="Paulmann" firstname="Clara Sophie" license="0">
              <RESULTS>
                <RESULT resultid="441" eventid="7" swimtime="00:01:25.60" reactiontime="+83" lane="5" heatid="7001" />
                <RESULT resultid="442" eventid="14" swimtime="00:00:40.80" lane="7" heatid="14002" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="162" birthdate="1998-01-01" gender="F" lastname="Gerungan" firstname="Daveena" license="0">
              <RESULTS>
                <RESULT resultid="443" eventid="7" swimtime="00:00:49.36" reactiontime="+92" lane="6" heatid="7008" />
                <RESULT resultid="444" eventid="14" swimtime="00:00:22.46" lane="7" heatid="14010" />
                <RESULT resultid="445" eventid="20" swimtime="00:01:52.92" reactiontime="+91" lane="7" heatid="20006">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:53.55" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="163" birthdate="2001-01-01" gender="M" lastname="Gaida" firstname="Duncan" license="0">
              <RESULTS>
                <RESULT resultid="446" eventid="2" swimtime="00:03:18.13" reactiontime="+98" lane="4" heatid="2004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:47.32" />
                    <SPLIT distance="200" swimtime="00:01:37.40" />
                    <SPLIT distance="300" swimtime="00:02:28.15" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="447" eventid="10" swimtime="00:06:46.45" reactiontime="+97" lane="4" heatid="10001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:47.16" />
                    <SPLIT distance="200" swimtime="00:01:37.36" />
                    <SPLIT distance="300" swimtime="00:02:28.59" />
                    <SPLIT distance="400" swimtime="00:03:20.66" />
                    <SPLIT distance="500" swimtime="00:04:12.78" />
                    <SPLIT distance="600" swimtime="00:05:05.30" />
                    <SPLIT distance="700" swimtime="00:05:57.06" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="164" birthdate="2007-01-01" gender="F" lastname="Hempler" firstname="Emily" license="0">
              <RESULTS>
                <RESULT resultid="448" eventid="1" status="DNS" swimtime="00:00:00.00" lane="3" heatid="1005" />
                <RESULT resultid="449" eventid="7" status="DNS" swimtime="00:00:00.00" lane="3" heatid="7009" />
                <RESULT resultid="450" eventid="14" status="DNS" swimtime="00:00:00.00" lane="4" heatid="14010" />
                <RESULT resultid="451" eventid="20" status="DNS" swimtime="00:00:00.00" lane="3" heatid="20007" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="165" birthdate="1999-01-01" gender="M" lastname="Wahlstadt" firstname="Felix" license="267">
              <RESULTS>
                <RESULT resultid="452" eventid="10" swimtime="00:07:26.98" reactiontime="+96" lane="3" heatid="10001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:49.35" />
                    <SPLIT distance="200" swimtime="00:01:43.32" />
                    <SPLIT distance="300" swimtime="00:02:38.94" />
                    <SPLIT distance="400" swimtime="00:03:35.44" />
                    <SPLIT distance="500" swimtime="00:04:32.67" />
                    <SPLIT distance="600" swimtime="00:05:30.34" />
                    <SPLIT distance="700" swimtime="00:06:28.93" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="453" eventid="15" swimtime="00:00:18.57" lane="3" heatid="15009" />
                <RESULT resultid="454" eventid="19" status="DNS" swimtime="00:00:00.00" lane="5" heatid="19002" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="166" birthdate="2011-01-01" gender="F" lastname="Hau" firstname="Hannah" license="0">
              <RESULTS>
                <RESULT resultid="455" eventid="7" swimtime="00:01:09.25" reactiontime="+73" lane="3" heatid="7003" />
                <RESULT resultid="456" eventid="14" swimtime="00:00:30.97" lane="5" heatid="14003" />
                <RESULT resultid="457" eventid="20" swimtime="00:02:33.41" lane="2" heatid="20003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:11.94" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="167" birthdate="2008-01-01" gender="F" lastname="Säbisch" firstname="Kyra" license="0">
              <RESULTS>
                <RESULT resultid="458" eventid="5" swimtime="00:00:20.86" lane="1" heatid="5003" />
                <RESULT resultid="459" eventid="7" swimtime="00:00:52.69" reactiontime="+97" lane="1" heatid="7008" />
                <RESULT resultid="460" eventid="20" swimtime="00:01:58.42" reactiontime="+96" lane="7" heatid="20005">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:55.45" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="168" birthdate="2008-01-01" gender="M" lastname="Hauk" firstname="Leon" license="0">
              <RESULTS>
                <RESULT resultid="461" eventid="6" swimtime="00:00:29.62" lane="3" heatid="6001" />
                <RESULT resultid="462" eventid="8" swimtime="00:01:11.66" reactiontime="+95" lane="3" heatid="8004" />
                <RESULT resultid="463" eventid="15" swimtime="00:00:30.58" lane="7" heatid="15005" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="169" birthdate="2007-01-01" gender="F" lastname="Holtz" firstname="Leonie-Florentine" license="2947">
              <RESULTS>
                <RESULT resultid="464" eventid="1" swimtime="00:04:28.80" reactiontime="+97" lane="1" heatid="1004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:00.21" />
                    <SPLIT distance="200" swimtime="00:02:09.64" />
                    <SPLIT distance="300" swimtime="00:03:20.10" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="465" eventid="14" swimtime="00:00:23.62" lane="2" heatid="14010" />
                <RESULT resultid="466" eventid="18" swimtime="00:00:52.99" reactiontime="+92" lane="2" heatid="18003" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="170" birthdate="2013-01-01" gender="F" lastname="Kannenberg" firstname="Lilly" license="0">
              <RESULTS>
                <RESULT resultid="467" eventid="7" swimtime="00:01:14.04" lane="5" heatid="7003" />
                <RESULT resultid="468" eventid="14" swimtime="00:00:32.79" lane="4" heatid="14003" />
                <RESULT resultid="469" eventid="20" swimtime="00:02:38.22" lane="8" heatid="20003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:18.04" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="171" birthdate="2008-01-01" gender="F" lastname="Horenok" firstname="Maiia" license="0">
              <RESULTS>
                <RESULT resultid="470" eventid="1" swimtime="00:03:41.92" reactiontime="+94" lane="2" heatid="1005">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:51.60" />
                    <SPLIT distance="200" swimtime="00:01:49.40" />
                    <SPLIT distance="300" swimtime="00:02:46.86" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="471" eventid="7" swimtime="00:00:44.90" reactiontime="+98" lane="3" heatid="7010" />
                <RESULT resultid="472" eventid="14" swimtime="00:00:19.68" lane="3" heatid="14011" />
                <RESULT resultid="473" eventid="18" swimtime="00:00:44.12" lane="5" heatid="18003" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="172" birthdate="2011-01-01" gender="F" lastname="Oesterreich" firstname="Mara" license="0">
              <RESULTS>
                <RESULT resultid="474" eventid="7" swimtime="00:01:16.37" lane="2" heatid="7002" />
                <RESULT resultid="475" eventid="14" swimtime="00:00:33.06" lane="5" heatid="14002" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="173" birthdate="2012-01-01" gender="M" lastname="Schnepel" firstname="Marten" license="0">
              <RESULTS>
                <RESULT resultid="476" eventid="8" status="DNS" swimtime="00:00:00.00" lane="5" heatid="8002" />
                <RESULT resultid="477" eventid="15" status="DNS" swimtime="00:00:00.00" lane="8" heatid="15003" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="174" birthdate="2011-01-01" gender="F" lastname="Schröter" firstname="Melissa" license="0">
              <RESULTS>
                <RESULT resultid="478" eventid="7" swimtime="00:01:15.07" lane="2" heatid="7003" />
                <RESULT resultid="479" eventid="14" swimtime="00:00:32.55" lane="1" heatid="14004" />
                <RESULT resultid="480" eventid="20" swimtime="00:02:49.67" lane="4" heatid="20002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:23.55" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="175" birthdate="2009-01-01" gender="M" lastname="Batiuk" firstname="Mykyta" license="0">
              <RESULTS>
                <RESULT resultid="481" eventid="6" swimtime="00:00:18.33" lane="8" heatid="6004" />
                <RESULT resultid="482" eventid="8" swimtime="00:00:46.35" reactiontime="+80" lane="4" heatid="8007" />
                <RESULT resultid="483" eventid="15" swimtime="00:00:20.57" lane="6" heatid="15008" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="176" birthdate="2012-01-01" gender="M" lastname="Kulchytskyi" firstname="Mykyta" license="0">
              <RESULTS>
                <RESULT resultid="484" eventid="8" swimtime="00:01:00.63" reactiontime="+96" lane="5" heatid="8004" />
                <RESULT resultid="485" eventid="15" swimtime="00:00:26.89" lane="5" heatid="15004" />
                <RESULT resultid="486" eventid="21" swimtime="00:02:16.59" reactiontime="+98" lane="6" heatid="21003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:04.35" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="177" birthdate="2004-01-01" gender="F" lastname="Barthel" firstname="Nadja" license="0">
              <RESULTS>
                <RESULT resultid="487" eventid="1" swimtime="00:03:46.59" reactiontime="+89" lane="3" heatid="1004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:50.62" />
                    <SPLIT distance="200" swimtime="00:01:48.46" />
                    <SPLIT distance="300" swimtime="00:02:48.16" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="488" eventid="5" swimtime="00:00:20.04" lane="1" heatid="5002" />
                <RESULT resultid="489" eventid="7" swimtime="00:00:45.64" reactiontime="+87" lane="8" heatid="7008" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="178" birthdate="2010-01-01" gender="F" lastname="Horenok" firstname="Polina" license="0">
              <RESULTS>
                <RESULT resultid="490" eventid="1" swimtime="00:04:43.88" reactiontime="+89" lane="2" heatid="1003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:05.33" />
                    <SPLIT distance="200" swimtime="00:02:20.45" />
                    <SPLIT distance="300" swimtime="00:03:36.00" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="491" eventid="7" swimtime="00:00:59.46" reactiontime="+91" lane="4" heatid="7006" />
                <RESULT resultid="492" eventid="14" swimtime="00:00:26.27" lane="6" heatid="14007" />
                <RESULT resultid="493" eventid="18" swimtime="00:01:05.41" lane="1" heatid="18002" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="179" birthdate="1998-01-01" gender="F" lastname="Niemann" firstname="Sophie" license="0">
              <RESULTS>
                <RESULT resultid="494" eventid="5" swimtime="00:00:18.56" lane="8" heatid="5004" />
                <RESULT resultid="495" eventid="7" swimtime="00:00:45.57" reactiontime="+94" lane="8" heatid="7010" />
                <RESULT resultid="496" eventid="14" swimtime="00:00:22.58" lane="7" heatid="14009" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="180" birthdate="2009-01-01" gender="F" lastname="Riekewald" firstname="Stella" license="0">
              <RESULTS>
                <RESULT resultid="497" eventid="5" swimtime="00:00:30.25" lane="8" heatid="5001" />
                <RESULT resultid="498" eventid="7" swimtime="00:01:17.30" lane="8" heatid="7004" />
                <RESULT resultid="499" eventid="14" swimtime="00:00:33.65" lane="7" heatid="14004" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="181" birthdate="2013-01-01" gender="F" lastname="Amelung" firstname="Tabea" license="0">
              <RESULTS>
                <RESULT resultid="500" eventid="7" status="DSQ" swimtime="00:00:41.45" reactiontime="+68" lane="1" heatid="7004" comment="Falscher Start." />
                <RESULT resultid="501" eventid="14" swimtime="00:00:30.57" lane="6" heatid="14004" />
                <RESULT resultid="502" eventid="20" swimtime="00:02:37.61" lane="7" heatid="20003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:18.67" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="184" birthdate="1976-01-01" gender="F" lastname="Paulmann" firstname="Anja" license="0">
              <RESULTS>
                <RESULT resultid="505" eventid="11" swimtime="00:00:27.82" lane="6" heatid="11001" />
                <RESULT resultid="506" eventid="14" swimtime="00:00:27.66" lane="6" heatid="14006" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="185" birthdate="1958-01-01" gender="F" lastname="Hirschfeldt" firstname="Birgit" license="0">
              <RESULTS>
                <RESULT resultid="507" eventid="11" swimtime="00:00:32.20" lane="2" heatid="11001" />
                <RESULT resultid="508" eventid="14" swimtime="00:00:30.86" lane="1" heatid="14006" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="186" birthdate="1987-01-01" gender="F" lastname="Eckstein" firstname="Diana" license="0">
              <RESULTS>
                <RESULT resultid="509" eventid="7" swimtime="00:00:57.18" reactiontime="+73" lane="2" heatid="7007" />
                <RESULT resultid="510" eventid="11" swimtime="00:00:27.58" lane="4" heatid="11001" />
                <RESULT resultid="511" eventid="14" swimtime="00:00:24.31" lane="2" heatid="14008" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="187" birthdate="1984-01-01" gender="F" lastname="Sapsai" firstname="Irina" license="0">
              <RESULTS>
                <RESULT resultid="512" eventid="11" swimtime="00:00:27.81" lane="3" heatid="11001" />
                <RESULT resultid="513" eventid="14" swimtime="00:00:28.17" lane="1" heatid="14008" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="188" birthdate="1978-01-01" gender="M" lastname="Bordag" firstname="Stefan" license="0">
              <RESULTS>
                <RESULT resultid="514" eventid="6" swimtime="00:00:22.58" lane="8" heatid="6003" />
                <RESULT resultid="515" eventid="8" swimtime="00:00:55.91" lane="6" heatid="8006" />
                <RESULT resultid="516" eventid="12" swimtime="00:00:26.60" lane="1" heatid="12002" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="189" birthdate="1977-01-01" gender="M" lastname="Nehrdich" firstname="Thomas" license="0">
              <RESULTS>
                <RESULT resultid="517" eventid="2" swimtime="00:03:55.46" reactiontime="+72" lane="4" heatid="2003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:51.99" />
                    <SPLIT distance="200" swimtime="00:01:52.57" />
                    <SPLIT distance="300" swimtime="00:02:56.13" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="518" eventid="8" swimtime="00:00:45.37" lane="3" heatid="8007" />
                <RESULT resultid="519" eventid="15" swimtime="00:00:19.84" lane="7" heatid="15008" />
                <RESULT resultid="520" eventid="21" swimtime="00:01:47.43" lane="4" heatid="21005">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:54.99" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="190" birthdate="1973-01-01" gender="M" lastname="Stelzig" firstname="Torsten" license="0">
              <RESULTS>
                <RESULT resultid="521" eventid="6" swimtime="00:00:22.37" lane="4" heatid="6002" />
                <RESULT resultid="522" eventid="12" swimtime="00:00:26.82" lane="4" heatid="12001" />
                <RESULT resultid="523" eventid="15" swimtime="00:00:24.73" lane="1" heatid="15007" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="191" birthdate="1969-01-01" gender="F" lastname="Meier-Mahlo" firstname="Ulrike" license="0">
              <RESULTS>
                <RESULT resultid="524" eventid="5" swimtime="00:00:22.42" lane="3" heatid="5002" />
                <RESULT resultid="525" eventid="11" swimtime="00:00:27.91" lane="5" heatid="11001" />
                <RESULT resultid="526" eventid="14" swimtime="00:00:24.36" lane="7" heatid="14008" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="192" birthdate="1967-01-01" gender="M" lastname="Meier" firstname="Wolf-Dieter" license="0">
              <RESULTS>
                <RESULT resultid="527" eventid="6" swimtime="00:00:20.89" lane="6" heatid="6003" />
                <RESULT resultid="528" eventid="8" swimtime="00:00:53.39" lane="7" heatid="8006" />
                <RESULT resultid="529" eventid="12" swimtime="00:00:25.47" lane="5" heatid="12002" />
                <RESULT resultid="530" eventid="15" swimtime="00:00:23.70" lane="6" heatid="15007" />
                <RESULT resultid="531" eventid="21" swimtime="00:02:05.20" lane="6" heatid="21005">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:59.58" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="290" birthdate="1987-01-01" gender="M" lastname="Eckstein" firstname="Diana" license="0" />
            <ATHLETE athleteid="294" birthdate="2008-01-01" gender="F" lastname="Kulchitska" firstname="Polina" license="0">
              <RESULTS>
                <RESULT resultid="706" eventid="1" swimtime="00:03:56.03" reactiontime="+93" lane="8" heatid="1005">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:54.74" />
                    <SPLIT distance="200" swimtime="00:01:56.42" />
                    <SPLIT distance="300" swimtime="00:02:57.20" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="707" eventid="9" swimtime="00:08:06.44" reactiontime="+93" lane="5" heatid="9002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:58.46" />
                    <SPLIT distance="200" swimtime="00:02:00.69" />
                    <SPLIT distance="300" swimtime="00:03:03.25" />
                    <SPLIT distance="400" swimtime="00:04:04.86" />
                    <SPLIT distance="500" swimtime="00:05:06.23" />
                    <SPLIT distance="600" swimtime="00:06:07.74" />
                    <SPLIT distance="700" swimtime="00:07:08.11" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="708" eventid="20" swimtime="00:01:53.16" lane="3" heatid="20006">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:54.75" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY number="1" gender="X" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="426" eventid="13" swimtime="00:01:22.33" lane="5" heatid="13002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:41.02" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="171" number="1" />
                    <RELAYPOSITION athleteid="158" number="2" />
                    <RELAYPOSITION athleteid="167" number="3" />
                    <RELAYPOSITION athleteid="160" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" gender="F" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="427" eventid="24" swimtime="00:03:17.86" lane="3" heatid="24002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:52.72" />
                    <SPLIT distance="200" swimtime="00:01:41.34" />
                    <SPLIT distance="300" swimtime="00:02:34.10" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="178" number="1" />
                    <RELAYPOSITION athleteid="162" number="2" />
                    <RELAYPOSITION athleteid="167" number="3" />
                    <RELAYPOSITION athleteid="171" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" gender="M" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="428" eventid="25" swimtime="00:02:48.75" lane="4" heatid="25001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:38.66" />
                    <SPLIT distance="200" swimtime="00:01:25.03" />
                    <SPLIT distance="300" swimtime="00:02:07.12" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="163" number="1" />
                    <RELAYPOSITION athleteid="158" number="2" />
                    <RELAYPOSITION athleteid="160" number="3" />
                    <RELAYPOSITION athleteid="165" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="2" gender="M" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="429" eventid="25" swimtime="00:04:41.64" lane="6" heatid="25001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:02.16" />
                    <SPLIT distance="200" swimtime="00:02:16.79" />
                    <SPLIT distance="300" swimtime="00:03:45.88" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="175" number="1" />
                    <RELAYPOSITION athleteid="168" number="2" />
                    <RELAYPOSITION athleteid="159" number="3" />
                    <RELAYPOSITION athleteid="173" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="2" gender="X" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="430" eventid="13" swimtime="00:02:01.66" lane="3" heatid="13001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:59.56" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="175" number="1" />
                    <RELAYPOSITION athleteid="180" number="2" />
                    <RELAYPOSITION athleteid="168" number="3" />
                    <RELAYPOSITION athleteid="166" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="2" gender="F" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="431" eventid="24" swimtime="00:04:47.32" lane="4" heatid="24001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:08.08" />
                    <SPLIT distance="200" swimtime="00:02:17.81" />
                    <SPLIT distance="300" swimtime="00:03:31.26" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="166" number="1" />
                    <RELAYPOSITION athleteid="181" number="2" />
                    <RELAYPOSITION athleteid="170" number="3" />
                    <RELAYPOSITION athleteid="174" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="3" gender="X" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="432" eventid="13" swimtime="00:02:25.61" lane="2" heatid="13001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:11.54" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="174" number="1" />
                    <RELAYPOSITION athleteid="159" number="2" />
                    <RELAYPOSITION athleteid="161" number="3" />
                    <RELAYPOSITION athleteid="172" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="100" gender="M" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="503" eventid="25" swimtime="00:03:44.05" lane="3" heatid="25001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:04.47" />
                    <SPLIT distance="200" swimtime="00:02:01.08" />
                    <SPLIT distance="300" swimtime="00:02:58.18" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="290" number="1" />
                    <RELAYPOSITION athleteid="190" number="2" />
                    <RELAYPOSITION athleteid="192" number="3" />
                    <RELAYPOSITION athleteid="189" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="100" gender="X" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="504" eventid="13" swimtime="00:01:40.91" lane="2" heatid="13002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:49.20" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="192" number="1" />
                    <RELAYPOSITION athleteid="187" number="2" />
                    <RELAYPOSITION athleteid="188" number="3" />
                    <RELAYPOSITION athleteid="191" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB name="SC Riesa Sekt. Flossenschwimmen" nation="GER" region="20" code="154149">
          <ATHLETES>
            <ATHLETE athleteid="141" birthdate="2011-01-01" gender="F" lastname="Hönisch" firstname="Ida" license="0">
              <RESULTS>
                <RESULT resultid="393" eventid="1" swimtime="00:05:19.30" reactiontime="+98" lane="5" heatid="1002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:10.11" />
                    <SPLIT distance="200" swimtime="00:02:31.90" />
                    <SPLIT distance="300" swimtime="00:03:56.19" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="394" eventid="7" swimtime="00:01:03.96" lane="5" heatid="7004" />
                <RESULT resultid="395" eventid="14" status="DSQ" swimtime="00:00:28.75" lane="3" heatid="14005" comment="Falscher Start." />
                <RESULT resultid="396" eventid="20" swimtime="00:02:24.22" lane="5" heatid="20003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:07.77" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="142" birthdate="2010-01-01" gender="F" lastname="Berger" firstname="Lene" license="0">
              <RESULTS>
                <RESULT resultid="397" eventid="1" swimtime="00:04:45.47" lane="4" heatid="1002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:05.16" />
                    <SPLIT distance="200" swimtime="00:02:17.44" />
                    <SPLIT distance="300" swimtime="00:03:33.00" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="398" eventid="7" swimtime="00:01:00.38" lane="4" heatid="7004" />
                <RESULT resultid="399" eventid="14" swimtime="00:00:27.63" lane="7" heatid="14006" />
                <RESULT resultid="400" eventid="20" swimtime="00:02:14.20" lane="2" heatid="20004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:04.61" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="143" birthdate="2014-01-01" gender="F" lastname="Näther" firstname="Mathilde" license="0">
              <RESULTS>
                <RESULT resultid="401" eventid="7" swimtime="00:01:50.00" reactiontime="+99" lane="6" heatid="7001" />
                <RESULT resultid="402" eventid="14" swimtime="00:00:49.90" lane="3" heatid="14001" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="144" birthdate="2014-01-01" gender="M" lastname="Fleck" firstname="Maximilian" license="0">
              <RESULTS>
                <RESULT resultid="403" eventid="8" swimtime="00:02:00.45" lane="6" heatid="8001" />
                <RESULT resultid="404" eventid="15" swimtime="00:00:53.08" lane="3" heatid="15001" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="146" birthdate="2014-01-01" gender="M" lastname="von Hoff" firstname="Neo" license="0">
              <RESULTS>
                <RESULT resultid="407" eventid="8" swimtime="00:01:42.60" reactiontime="+77" lane="5" heatid="8001" />
                <RESULT resultid="408" eventid="15" swimtime="00:00:43.75" lane="5" heatid="15001" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="147" birthdate="2006-01-01" gender="M" lastname="Loßner" firstname="Niklas" license="0">
              <RESULTS>
                <RESULT resultid="409" eventid="2" swimtime="00:03:37.87" reactiontime="+98" lane="3" heatid="2004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:48.44" />
                    <SPLIT distance="200" swimtime="00:01:45.03" />
                    <SPLIT distance="300" swimtime="00:02:43.02" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="410" eventid="8" swimtime="00:00:38.10" reactiontime="+93" lane="5" heatid="8008" />
                <RESULT resultid="411" eventid="15" swimtime="00:00:16.56" lane="5" heatid="15009" />
                <RESULT resultid="412" eventid="21" swimtime="00:01:37.42" reactiontime="+97" lane="3" heatid="21006">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:46.27" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="SG Dresden" nation="GER" region="20" code="0">
          <ATHLETES>
            <ATHLETE athleteid="263" birthdate="2012-01-01" gender="F" lastname="Bernhardt" firstname="Fjora" license="0">
              <RESULTS>
                <RESULT resultid="583" eventid="7" swimtime="00:01:16.88" lane="6" heatid="7003" />
                <RESULT resultid="584" eventid="14" swimtime="00:00:34.59" lane="3" heatid="14003" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="264" birthdate="1987-01-01" gender="M" lastname="Böhme" firstname="Johannes" license="0">
              <RESULTS>
                <RESULT resultid="585" eventid="2" swimtime="00:03:48.07" reactiontime="+90" lane="7" heatid="2004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:50.40" />
                    <SPLIT distance="200" swimtime="00:01:48.18" />
                    <SPLIT distance="300" swimtime="00:02:48.07" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="586" eventid="8" swimtime="00:00:46.96" reactiontime="+90" lane="5" heatid="8007" />
                <RESULT resultid="587" eventid="21" swimtime="00:01:44.81" reactiontime="+93" lane="8" heatid="21006">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:49.64" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="265" birthdate="2007-01-01" gender="F" lastname="Bretschneider" firstname="Luisa" license="0">
              <RESULTS>
                <RESULT resultid="588" eventid="5" swimtime="00:00:28.94" lane="7" heatid="5001" />
                <RESULT resultid="589" eventid="7" swimtime="00:01:10.74" reactiontime="+95" lane="3" heatid="7004" />
                <RESULT resultid="590" eventid="14" swimtime="00:00:30.50" lane="7" heatid="14005" />
                <RESULT resultid="591" eventid="20" swimtime="00:02:37.63" lane="6" heatid="20003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:14.63" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="266" birthdate="2011-01-01" gender="M" lastname="Buchmann" firstname="Marco" license="0">
              <RESULTS>
                <RESULT resultid="592" eventid="8" status="DNS" swimtime="00:00:00.00" lane="8" heatid="8004" />
                <RESULT resultid="593" eventid="15" status="DNS" swimtime="00:00:00.00" lane="4" heatid="15004" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="268" birthdate="1978-01-01" gender="M" lastname="Hoffmann" firstname="Stefan" license="0">
              <RESULTS>
                <RESULT resultid="598" eventid="6" swimtime="00:00:19.05" lane="7" heatid="6003" />
                <RESULT resultid="599" eventid="12" swimtime="00:00:23.39" lane="6" heatid="12002" />
                <RESULT resultid="600" eventid="15" swimtime="00:00:22.97" lane="2" heatid="15007" />
                <RESULT resultid="601" eventid="19" swimtime="00:00:47.75" reactiontime="+99" lane="5" heatid="19001" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="269" birthdate="2009-01-01" gender="M" lastname="Hübner" firstname="Christoph" license="0">
              <RESULTS>
                <RESULT resultid="602" eventid="8" swimtime="00:01:15.74" reactiontime="+99" lane="8" heatid="8003" />
                <RESULT resultid="603" eventid="15" swimtime="00:00:31.57" lane="5" heatid="15003" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="270" birthdate="1986-01-01" gender="F" lastname="Klar" firstname="Margarethe" license="0">
              <RESULTS>
                <RESULT resultid="604" eventid="1" swimtime="00:04:36.23" lane="5" heatid="1003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:02.65" />
                    <SPLIT distance="200" swimtime="00:02:13.95" />
                    <SPLIT distance="300" swimtime="00:03:26.27" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="605" eventid="7" swimtime="00:01:00.21" reactiontime="+98" lane="8" heatid="7007" />
                <RESULT resultid="606" eventid="14" swimtime="00:00:27.93" lane="4" heatid="14006" />
                <RESULT resultid="607" eventid="18" swimtime="00:00:59.15" lane="4" heatid="18002" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="271" birthdate="2009-01-01" gender="M" lastname="Lange" firstname="Viktor" license="0">
              <RESULTS>
                <RESULT resultid="608" eventid="8" swimtime="00:01:15.12" reactiontime="+97" lane="1" heatid="8003" />
                <RESULT resultid="609" eventid="15" swimtime="00:00:33.63" lane="3" heatid="15003" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="272" birthdate="2007-01-01" gender="F" lastname="Marquardt" firstname="Lotte" license="0">
              <RESULTS>
                <RESULT resultid="610" eventid="5" swimtime="00:00:25.79" lane="7" heatid="5002" />
                <RESULT resultid="611" eventid="7" swimtime="00:01:00.20" lane="1" heatid="7006" />
                <RESULT resultid="612" eventid="14" swimtime="00:00:27.98" lane="7" heatid="14007" />
                <RESULT resultid="613" eventid="18" swimtime="00:01:06.68" lane="8" heatid="18002" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="273" birthdate="2010-01-01" gender="F" lastname="Mucha" firstname="Helene" license="0">
              <RESULTS>
                <RESULT resultid="614" eventid="7" status="DSQ" swimtime="00:00:22.31" reactiontime="+87" lane="2" heatid="7004" comment="Aufgegeben nach 5 Meter." />
                <RESULT resultid="615" eventid="14" swimtime="00:00:32.42" lane="8" heatid="14005" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="274" birthdate="2011-01-01" gender="F" lastname="Müller" firstname="Reni" license="0">
              <RESULTS>
                <RESULT resultid="616" eventid="7" swimtime="00:01:13.36" reactiontime="+81" lane="7" heatid="7004" />
                <RESULT resultid="617" eventid="14" swimtime="00:00:31.03" lane="4" heatid="14004" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="275" birthdate="2006-01-01" gender="F" lastname="Neumann" firstname="Josephine" license="0">
              <RESULTS>
                <RESULT resultid="618" eventid="5" swimtime="00:00:26.32" lane="3" heatid="5001" />
                <RESULT resultid="619" eventid="7" swimtime="00:01:01.92" reactiontime="+98" lane="7" heatid="7006" />
                <RESULT resultid="620" eventid="14" swimtime="00:00:28.21" lane="5" heatid="14006" />
                <RESULT resultid="621" eventid="20" swimtime="00:02:21.24" reactiontime="+98" lane="8" heatid="20005">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:08.06" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="276" birthdate="2011-01-01" gender="F" lastname="Oehme" firstname="Mia" license="0">
              <RESULTS>
                <RESULT resultid="622" eventid="7" swimtime="00:01:10.98" reactiontime="+95" lane="8" heatid="7003" />
                <RESULT resultid="623" eventid="14" swimtime="00:00:31.57" lane="8" heatid="14004" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="277" birthdate="1999-01-01" gender="M" lastname="Petrich" firstname="Mike" license="0">
              <RESULTS>
                <RESULT resultid="624" eventid="23" swimtime="00:04:46.11" lane="2" heatid="23001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:01.34" />
                    <SPLIT distance="200" swimtime="00:02:15.30" />
                    <SPLIT distance="300" swimtime="00:03:32.19" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="278" birthdate="2005-01-01" gender="M" lastname="Petrich" firstname="Nick" license="0">
              <RESULTS>
                <RESULT resultid="625" eventid="23" status="DSQ" swimtime="00:05:54.59" lane="7" heatid="23001" comment="Falsche Wende bei 100m.">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:15.70" />
                    <SPLIT distance="200" swimtime="00:02:50.72" />
                    <SPLIT distance="300" swimtime="00:04:24.41" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="279" birthdate="2004-01-01" gender="F" lastname="Placzek" firstname="Lilly" license="0">
              <RESULTS>
                <RESULT resultid="626" eventid="5" swimtime="00:00:17.91" lane="3" heatid="5004" />
                <RESULT resultid="627" eventid="7" swimtime="00:00:46.63" reactiontime="+95" lane="7" heatid="7010" />
                <RESULT resultid="628" eventid="14" swimtime="00:00:20.13" lane="6" heatid="14011" />
                <RESULT resultid="629" eventid="18" swimtime="00:00:44.58" reactiontime="+90" lane="5" heatid="18004" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="280" birthdate="2007-01-01" gender="F" lastname="Razumovska" firstname="Sophia" license="0">
              <RESULTS>
                <RESULT resultid="630" eventid="5" swimtime="00:00:28.16" lane="2" heatid="5001" />
                <RESULT resultid="631" eventid="7" swimtime="00:01:05.94" reactiontime="+90" lane="3" heatid="7005" />
                <RESULT resultid="632" eventid="14" swimtime="00:00:29.01" lane="2" heatid="14006" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="281" birthdate="2010-01-01" gender="F" lastname="Reichel" firstname="Emily" license="0">
              <RESULTS>
                <RESULT resultid="633" eventid="7" swimtime="00:01:05.24" reactiontime="+99" lane="1" heatid="7005" />
                <RESULT resultid="634" eventid="14" swimtime="00:00:28.65" lane="8" heatid="14006" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="282" birthdate="2005-01-01" gender="F" lastname="Richter" firstname="Franca" license="0">
              <RESULTS>
                <RESULT resultid="635" eventid="1" swimtime="00:03:51.95" reactiontime="+99" lane="5" heatid="1005">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:53.78" />
                    <SPLIT distance="200" swimtime="00:01:52.97" />
                    <SPLIT distance="300" swimtime="00:02:52.55" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="636" eventid="18" swimtime="00:00:41.68" lane="3" heatid="18004" />
                <RESULT resultid="637" eventid="20" swimtime="00:01:42.28" lane="7" heatid="20007">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:49.46" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="283" birthdate="2000-01-01" gender="F" lastname="Rütze" firstname="Michele" license="0">
              <RESULTS>
                <RESULT resultid="639" eventid="5" swimtime="00:00:17.11" lane="4" heatid="5004" />
                <RESULT resultid="640" eventid="7" swimtime="00:00:40.98" reactiontime="+87" lane="4" heatid="7010" />
                <RESULT resultid="641" eventid="14" swimtime="00:00:18.99" lane="4" heatid="14011" />
                <RESULT resultid="642" eventid="18" swimtime="00:00:39.73" lane="4" heatid="18004" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="284" birthdate="2006-01-01" gender="F" lastname="Schürer" firstname="Katka" license="0">
              <RESULTS>
                <RESULT resultid="643" eventid="7" status="DSQ" swimtime="00:01:10.99" reactiontime="+59" lane="7" heatid="7003" comment="Falscher Start." />
                <RESULT resultid="644" eventid="14" swimtime="00:00:30.66" lane="6" heatid="14003" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="288" birthdate="2013-01-01" gender="F" lastname="Stegmann" firstname="Anna" license="0">
              <RESULTS>
                <RESULT resultid="648" eventid="7" status="DSQ" swimtime="00:01:16.20" lane="4" heatid="7002" comment="Falscher Start." />
                <RESULT resultid="649" eventid="14" swimtime="00:00:32.55" lane="8" heatid="14003" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="289" birthdate="2005-01-01" gender="F" lastname="Wielens" firstname="Hellen" license="0">
              <RESULTS>
                <RESULT resultid="650" eventid="22" swimtime="00:06:04.90" lane="1" heatid="22001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:23.89" />
                    <SPLIT distance="200" swimtime="00:02:55.85" />
                    <SPLIT distance="300" swimtime="00:04:28.68" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="291" birthdate="2002-01-01" gender="F" lastname="Klabunde" firstname="Lotte" license="0">
              <RESULTS>
                <RESULT resultid="652" eventid="1" swimtime="00:03:47.49" reactiontime="+97" lane="6" heatid="1004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:53.99" />
                    <SPLIT distance="200" swimtime="00:01:51.55" />
                    <SPLIT distance="300" swimtime="00:02:50.88" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="654" eventid="5" swimtime="00:00:19.99" lane="2" heatid="5004" />
                <RESULT resultid="653" eventid="7" status="WDR" swimtime="00:00:00.00" lane="2" heatid="7001" />
                <RESULT resultid="721" eventid="9" swimtime="00:08:26.34" reactiontime="+99" lane="6" heatid="9001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:57.90" />
                    <SPLIT distance="200" swimtime="00:02:00.53" />
                    <SPLIT distance="300" swimtime="00:03:04.60" />
                    <SPLIT distance="400" swimtime="00:04:09.08" />
                    <SPLIT distance="500" swimtime="00:05:13.95" />
                    <SPLIT distance="600" swimtime="00:06:20.40" />
                    <SPLIT distance="700" swimtime="00:07:27.40" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="655" eventid="18" swimtime="00:00:46.52" lane="2" heatid="18004" />
                <RESULT resultid="656" eventid="20" swimtime="00:01:46.48" reactiontime="+99" lane="8" heatid="20007">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:51.84" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="657" eventid="22" swimtime="00:04:03.91" lane="3" heatid="22001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:52.84" />
                    <SPLIT distance="200" swimtime="00:01:54.59" />
                    <SPLIT distance="300" swimtime="00:03:01.05" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY number="1" gender="F" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="645" eventid="24" status="DSQ" swimtime="00:03:01.66" lane="5" heatid="24002" comment="2. Starter: 15m nach dem Start übertaucht.">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:45.51" />
                    <SPLIT distance="200" swimtime="00:01:31.85" />
                    <SPLIT distance="300" swimtime="00:02:20.34" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="282" number="1" />
                    <RELAYPOSITION athleteid="279" number="2" />
                    <RELAYPOSITION athleteid="291" number="3" />
                    <RELAYPOSITION athleteid="283" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="2" gender="F" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="646" eventid="24" swimtime="00:04:24.23" lane="1" heatid="24002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:02.74" />
                    <SPLIT distance="200" swimtime="00:02:10.22" />
                    <SPLIT distance="300" swimtime="00:03:20.94" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="272" number="1" />
                    <RELAYPOSITION athleteid="280" number="2" />
                    <RELAYPOSITION athleteid="265" number="3" />
                    <RELAYPOSITION athleteid="275" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="3" gender="F" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="647" eventid="24" swimtime="00:04:58.03" lane="5" heatid="24001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:16.39" />
                    <SPLIT distance="200" swimtime="00:02:27.89" />
                    <SPLIT distance="300" swimtime="00:03:47.53" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="273" number="1" />
                    <RELAYPOSITION athleteid="276" number="2" />
                    <RELAYPOSITION athleteid="288" number="3" />
                    <RELAYPOSITION athleteid="274" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB name="SSC Halle" nation="GER" region="27" code="0">
          <ATHLETES>
            <ATHLETE athleteid="82" birthdate="2007-01-01" gender="M" lastname="Koch" firstname="Elias" license="0">
              <RESULTS>
                <RESULT resultid="215" eventid="6" swimtime="00:00:19.45" lane="4" heatid="6003" />
                <RESULT resultid="216" eventid="8" status="DSQ" swimtime="00:00:48.20" reactiontime="+88" lane="6" heatid="8007" comment="15m nach Start übertaucht." />
                <RESULT resultid="217" eventid="15" status="DSQ" swimtime="00:00:21.81" lane="4" heatid="15007" comment="15m nach Start übertaucht." />
                <RESULT resultid="218" eventid="19" swimtime="00:00:53.19" lane="1" heatid="19002" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="83" birthdate="2010-01-01" gender="M" lastname="Eichberg" firstname="Eric" license="0">
              <RESULTS>
                <RESULT resultid="219" eventid="8" status="DSQ" swimtime="00:01:15.27" lane="4" heatid="8002" comment="15m nach Start übertaucht." />
                <RESULT resultid="220" eventid="15" swimtime="00:00:37.74" lane="6" heatid="15003" />
                <RESULT resultid="221" eventid="21" swimtime="00:02:47.17" reactiontime="+86" lane="8" heatid="21003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:22.59" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="84" birthdate="2008-01-01" gender="M" lastname="Baumbach" firstname="Felix" license="0">
              <RESULTS>
                <RESULT resultid="222" eventid="2" status="DNS" swimtime="00:00:00.00" lane="3" heatid="2003" />
                <RESULT resultid="223" eventid="8" status="DNS" swimtime="00:00:00.00" lane="7" heatid="8007" />
                <RESULT resultid="224" eventid="10" status="WDR" swimtime="00:00:00.00" lane="0" heatid="10000" />
                <RESULT resultid="225" eventid="21" status="DNS" swimtime="00:00:00.00" lane="5" heatid="21005" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="85" birthdate="2013-01-01" gender="M" lastname="Rosemann" firstname="Henri" license="0">
              <RESULTS>
                <RESULT resultid="226" eventid="8" swimtime="00:01:15.77" reactiontime="+99" lane="3" heatid="8003" />
                <RESULT resultid="227" eventid="15" swimtime="00:00:35.37" lane="7" heatid="15003" />
                <RESULT resultid="228" eventid="21" status="DSQ" swimtime="00:00:00.00" lane="7" heatid="21002" comment="Aufgegeben nach 110 Meter.">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:24.17" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="86" birthdate="2011-01-01" gender="M" lastname="Reinicke" firstname="Jakob" license="0">
              <RESULTS>
                <RESULT resultid="229" eventid="2" swimtime="00:05:14.54" reactiontime="+73" lane="5" heatid="2002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:13.95" />
                    <SPLIT distance="200" swimtime="00:02:36.45" />
                    <SPLIT distance="300" swimtime="00:03:58.89" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="230" eventid="8" swimtime="00:01:01.54" reactiontime="+81" lane="6" heatid="8005" />
                <RESULT resultid="231" eventid="15" swimtime="00:00:27.51" lane="2" heatid="15006" />
                <RESULT resultid="232" eventid="21" swimtime="00:02:12.26" reactiontime="+87" lane="5" heatid="21003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:03.21" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="87" birthdate="2010-01-01" gender="M" lastname="Harms" firstname="Justus" license="0">
              <RESULTS>
                <RESULT resultid="233" eventid="2" swimtime="00:05:54.99" reactiontime="+78" lane="1" heatid="2003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:20.17" />
                    <SPLIT distance="200" swimtime="00:02:54.85" />
                    <SPLIT distance="300" swimtime="00:04:29.86" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="234" eventid="8" swimtime="00:01:02.72" reactiontime="+74" lane="3" heatid="8005" />
                <RESULT resultid="235" eventid="15" swimtime="00:00:27.76" lane="8" heatid="15006" />
                <RESULT resultid="236" eventid="21" swimtime="00:02:31.83" reactiontime="+78" lane="1" heatid="21004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:14.56" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="88" birthdate="2007-01-01" gender="F" lastname="Gallitz" firstname="Laura" license="0">
              <RESULTS>
                <RESULT resultid="237" eventid="5" swimtime="00:00:24.48" lane="4" heatid="5001" />
                <RESULT resultid="238" eventid="7" status="DSQ" swimtime="00:00:58.45" lane="1" heatid="7007" comment="15m nach Start übertaucht." />
                <RESULT resultid="239" eventid="14" swimtime="00:00:25.70" lane="2" heatid="14007" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="89" birthdate="2006-01-01" gender="F" lastname="Dietrich" firstname="Lea" license="0">
              <RESULTS>
                <RESULT resultid="240" eventid="5" swimtime="00:00:20.68" lane="5" heatid="5003" />
                <RESULT resultid="241" eventid="7" swimtime="00:00:49.55" reactiontime="+95" lane="8" heatid="7009" />
                <RESULT resultid="242" eventid="14" swimtime="00:00:21.98" lane="1" heatid="14010" />
                <RESULT resultid="243" eventid="20" swimtime="00:01:55.21" reactiontime="+94" lane="2" heatid="20006">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:55.04" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="90" birthdate="2013-01-01" gender="F" lastname="Wilke" firstname="Lieselotte" license="0">
              <RESULTS>
                <RESULT resultid="244" eventid="7" swimtime="00:01:22.33" reactiontime="+89" lane="1" heatid="7003" />
                <RESULT resultid="245" eventid="14" swimtime="00:00:36.97" lane="1" heatid="14003" />
                <RESULT resultid="246" eventid="20" status="DNS" swimtime="00:00:00.00" lane="5" heatid="20002" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="91" birthdate="2013-01-01" gender="F" lastname="Wilke" firstname="Martha" license="0">
              <RESULTS>
                <RESULT resultid="247" eventid="7" swimtime="00:01:15.50" reactiontime="+96" lane="7" heatid="7002" />
                <RESULT resultid="248" eventid="14" swimtime="00:00:33.24" lane="6" heatid="14002" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="93" birthdate="2007-01-01" gender="F" lastname="Gerlach" firstname="Meret" license="0">
              <RESULTS>
                <RESULT resultid="251" eventid="1" swimtime="00:04:10.55" reactiontime="+90" lane="2" heatid="1004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:58.50" />
                    <SPLIT distance="200" swimtime="00:02:03.23" />
                    <SPLIT distance="300" swimtime="00:03:06.82" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="252" eventid="9" swimtime="00:08:35.48" lane="6" heatid="9002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:59.74" />
                    <SPLIT distance="200" swimtime="00:02:04.29" />
                    <SPLIT distance="300" swimtime="00:03:09.81" />
                    <SPLIT distance="400" swimtime="00:04:15.41" />
                    <SPLIT distance="500" swimtime="00:05:21.83" />
                    <SPLIT distance="600" swimtime="00:06:28.62" />
                    <SPLIT distance="700" swimtime="00:07:33.53" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="253" eventid="14" swimtime="00:00:23.72" lane="2" heatid="14009" />
                <RESULT resultid="254" eventid="20" swimtime="00:01:56.97" reactiontime="+96" lane="6" heatid="20006">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:56.81" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="94" birthdate="2009-01-01" gender="M" lastname="Gaudig" firstname="Paul" license="0">
              <RESULTS>
                <RESULT resultid="255" eventid="6" swimtime="00:00:23.84" lane="7" heatid="6002" />
                <RESULT resultid="256" eventid="8" swimtime="00:00:54.53" lane="1" heatid="8005" />
                <RESULT resultid="257" eventid="15" swimtime="00:00:24.35" lane="6" heatid="15006" />
                <RESULT resultid="258" eventid="21" swimtime="00:02:12.77" lane="2" heatid="21004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:01.86" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="95" birthdate="2011-01-01" gender="M" lastname="Frenzel" firstname="Tim" license="0">
              <RESULTS>
                <RESULT resultid="259" eventid="2" swimtime="00:05:28.84" reactiontime="+96" lane="3" heatid="2002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:16.18" />
                    <SPLIT distance="200" swimtime="00:02:40.83" />
                    <SPLIT distance="300" swimtime="00:04:09.36" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="260" eventid="8" swimtime="00:01:11.10" lane="6" heatid="8004" />
                <RESULT resultid="261" eventid="15" swimtime="00:00:29.97" lane="8" heatid="15005" />
                <RESULT resultid="262" eventid="21" swimtime="00:02:39.32" lane="2" heatid="21003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:17.17" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="96" birthdate="2012-01-01" gender="M" lastname="Gaudig" firstname="Tom" license="0">
              <RESULTS>
                <RESULT resultid="263" eventid="8" swimtime="00:01:11.35" lane="4" heatid="8003" />
                <RESULT resultid="264" eventid="15" swimtime="00:00:32.95" lane="6" heatid="15004" />
                <RESULT resultid="265" eventid="21" swimtime="00:02:47.62" reactiontime="+95" lane="7" heatid="21003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:22.11" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY number="1" gender="X" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="266" eventid="13" swimtime="00:01:29.93" lane="3" heatid="13002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:46.00" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="89" number="1" />
                    <RELAYPOSITION athleteid="94" number="2" />
                    <RELAYPOSITION athleteid="82" number="3" />
                    <RELAYPOSITION athleteid="93" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="2" gender="X" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="267" eventid="13" swimtime="00:02:19.22" lane="5" heatid="13001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:06.54" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="96" number="1" />
                    <RELAYPOSITION athleteid="91" number="2" />
                    <RELAYPOSITION athleteid="85" number="3" />
                    <RELAYPOSITION athleteid="90" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB name="Tauchclub Jena" nation="GER" region="35" code="0">
          <ATHLETES>
            <ATHLETE athleteid="6" birthdate="2008-01-01" gender="M" lastname="Steininger" firstname="Bruno" license="0">
              <RESULTS>
                <RESULT resultid="23" eventid="2" swimtime="00:04:19.78" lane="5" heatid="2003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:00.56" />
                    <SPLIT distance="200" swimtime="00:02:06.11" />
                    <SPLIT distance="300" swimtime="00:03:14.37" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="24" eventid="6" status="DSQ" swimtime="00:00:00.00" lane="5" heatid="6002" comment="Gesicht aus dem Wasser bei 10 Meter." />
                <RESULT resultid="25" eventid="19" swimtime="00:00:52.20" lane="3" heatid="19001" />
                <RESULT resultid="26" eventid="21" swimtime="00:01:57.08" lane="3" heatid="21005">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:56.89" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="7" birthdate="1999-01-01" gender="F" lastname="Jacke" firstname="Lena" license="0">
              <RESULTS>
                <RESULT resultid="27" eventid="1" swimtime="00:04:12.32" reactiontime="+97" lane="7" heatid="1004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:02.27" />
                    <SPLIT distance="200" swimtime="00:02:06.62" />
                    <SPLIT distance="300" swimtime="00:03:11.80" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="28" eventid="9" swimtime="00:08:51.61" lane="2" heatid="9002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:04.51" />
                    <SPLIT distance="200" swimtime="00:02:09.88" />
                    <SPLIT distance="300" swimtime="00:03:15.09" />
                    <SPLIT distance="400" swimtime="00:04:24.75" />
                    <SPLIT distance="500" swimtime="00:05:31.70" />
                    <SPLIT distance="600" swimtime="00:06:38.09" />
                    <SPLIT distance="700" swimtime="00:07:48.87" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="29" eventid="16" swimtime="00:16:57.23" reactiontime="+98" lane="5" heatid="16001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:03.75" />
                    <SPLIT distance="200" swimtime="00:02:09.41" />
                    <SPLIT distance="300" swimtime="00:03:20.37" />
                    <SPLIT distance="400" swimtime="00:04:26.58" />
                    <SPLIT distance="500" swimtime="00:05:37.76" />
                    <SPLIT distance="600" swimtime="00:06:44.33" />
                    <SPLIT distance="700" swimtime="00:07:57.21" />
                    <SPLIT distance="800" swimtime="00:09:03.49" />
                    <SPLIT distance="900" swimtime="00:10:15.07" />
                    <SPLIT distance="1000" swimtime="00:11:20.65" />
                    <SPLIT distance="1100" swimtime="00:12:31.78" />
                    <SPLIT distance="1200" swimtime="00:13:37.75" />
                    <SPLIT distance="1300" swimtime="00:14:48.27" />
                    <SPLIT distance="1400" swimtime="00:15:55.47" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="30" eventid="22" swimtime="00:04:23.89" lane="7" heatid="22001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:00.74" />
                    <SPLIT distance="200" swimtime="00:02:05.75" />
                    <SPLIT distance="300" swimtime="00:03:17.69" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="8" birthdate="2009-01-01" gender="F" lastname="Steininger" firstname="Magda" license="0">
              <RESULTS>
                <RESULT resultid="31" eventid="5" swimtime="00:00:24.66" lane="8" heatid="5002" />
                <RESULT resultid="32" eventid="7" swimtime="00:00:57.74" reactiontime="+98" lane="3" heatid="7006" />
                <RESULT resultid="33" eventid="18" swimtime="00:00:58.98" lane="6" heatid="18002" />
                <RESULT resultid="34" eventid="20" swimtime="00:02:08.28" reactiontime="+77" lane="1" heatid="20005">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:01.54" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="9" birthdate="2005-01-01" gender="M" lastname="Preuß" firstname="Marek" license="0">
              <RESULTS>
                <RESULT resultid="35" eventid="2" swimtime="00:03:45.04" reactiontime="+79" lane="8" heatid="2004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:56.41" />
                    <SPLIT distance="200" swimtime="00:01:54.04" />
                    <SPLIT distance="300" swimtime="00:02:48.67" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="36" eventid="10" swimtime="00:08:04.54" reactiontime="+82" lane="2" heatid="10001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:59.18" />
                    <SPLIT distance="200" swimtime="00:01:59.62" />
                    <SPLIT distance="300" swimtime="00:02:57.15" />
                    <SPLIT distance="400" swimtime="00:04:02.19" />
                    <SPLIT distance="500" swimtime="00:05:04.65" />
                    <SPLIT distance="600" swimtime="00:06:03.54" />
                    <SPLIT distance="700" swimtime="00:07:08.74" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="37" eventid="19" swimtime="00:00:43.42" lane="7" heatid="19002" />
                <RESULT resultid="38" eventid="23" swimtime="00:03:39.40" lane="6" heatid="23001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:50.23" />
                    <SPLIT distance="200" swimtime="00:01:45.01" />
                    <SPLIT distance="300" swimtime="00:02:44.72" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="Tauchclub NEMO Plauen e.V." nation="GER" region="20" code="0">
          <ATHLETES>
            <ATHLETE athleteid="121" birthdate="1955-01-01" gender="M" lastname="Reuter" firstname="Andreas" license="0">
              <RESULTS>
                <RESULT resultid="324" eventid="6" swimtime="00:00:25.93" lane="2" heatid="6002" />
                <RESULT resultid="325" eventid="8" swimtime="00:01:05.36" lane="8" heatid="8005" />
                <RESULT resultid="326" eventid="12" swimtime="00:00:29.94" lane="3" heatid="12001" />
                <RESULT resultid="327" eventid="15" swimtime="00:00:29.01" lane="1" heatid="15006" />
                <RESULT resultid="328" eventid="19" swimtime="00:01:01.96" lane="2" heatid="19001" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="122" birthdate="2013-01-01" gender="M" lastname="Hertel" firstname="Etienne" license="0">
              <RESULTS>
                <RESULT resultid="329" eventid="2" swimtime="00:06:39.82" lane="3" heatid="2001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:33.05" />
                    <SPLIT distance="200" swimtime="00:03:17.43" />
                    <SPLIT distance="300" swimtime="00:05:00.22" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="330" eventid="8" swimtime="00:01:31.59" lane="7" heatid="8002" />
                <RESULT resultid="331" eventid="15" swimtime="00:00:40.14" lane="3" heatid="15002" />
                <RESULT resultid="332" eventid="21" swimtime="00:03:16.69" reactiontime="+84" lane="6" heatid="21001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:34.76" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="123" birthdate="2009-01-01" gender="F" lastname="Troppschuh" firstname="Hannah" license="0">
              <RESULTS>
                <RESULT resultid="333" eventid="5" swimtime="00:00:19.03" lane="7" heatid="5004" />
                <RESULT resultid="334" eventid="7" swimtime="00:00:46.44" reactiontime="+96" lane="4" heatid="7009" />
                <RESULT resultid="335" eventid="14" swimtime="00:00:22.07" lane="6" heatid="14010" />
                <RESULT resultid="336" eventid="18" swimtime="00:00:45.27" lane="7" heatid="18004" />
                <RESULT resultid="705" eventid="22" swimtime="00:03:44.22" lane="4" heatid="22001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:49.31" />
                    <SPLIT distance="200" swimtime="00:01:45.94" />
                    <SPLIT distance="300" swimtime="00:02:45.86" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="124" birthdate="2003-01-01" gender="F" lastname="Prochaska" firstname="Julia" license="0">
              <RESULTS>
                <RESULT resultid="338" eventid="5" swimtime="00:00:20.65" lane="7" heatid="5003" />
                <RESULT resultid="339" eventid="7" swimtime="00:00:52.24" lane="1" heatid="7009" />
                <RESULT resultid="340" eventid="14" swimtime="00:00:23.12" lane="4" heatid="14009" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="125" birthdate="2010-01-01" gender="F" lastname="Dawert" firstname="Klara" license="0">
              <RESULTS>
                <RESULT resultid="341" eventid="7" swimtime="00:01:13.57" lane="8" heatid="7005" />
                <RESULT resultid="342" eventid="14" swimtime="00:00:33.11" lane="1" heatid="14005" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="126" birthdate="2013-01-01" gender="F" lastname="Küthemann" firstname="Lina" license="0">
              <RESULTS>
                <RESULT resultid="343" eventid="1" status="WDR" swimtime="00:00:00.00" lane="3" heatid="1001" />
                <RESULT resultid="344" eventid="7" status="WDR" swimtime="00:00:00.00" lane="6" heatid="7002" />
                <RESULT resultid="345" eventid="14" status="WDR" swimtime="00:00:00.00" lane="2" heatid="14003" />
                <RESULT resultid="346" eventid="20" status="WDR" swimtime="00:00:00.00" lane="7" heatid="20002" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="127" birthdate="2012-01-01" gender="F" lastname="Troppschuh" firstname="Lotte" license="0">
              <RESULTS>
                <RESULT resultid="347" eventid="1" swimtime="00:04:45.17" reactiontime="+92" lane="6" heatid="1003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:05.67" />
                    <SPLIT distance="200" swimtime="00:02:18.88" />
                    <SPLIT distance="300" swimtime="00:03:32.91" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="348" eventid="7" swimtime="00:00:53.82" reactiontime="+94" lane="4" heatid="7007" />
                <RESULT resultid="349" eventid="14" swimtime="00:00:23.28" lane="4" heatid="14008" />
                <RESULT resultid="350" eventid="20" swimtime="00:02:10.04" reactiontime="+98" lane="6" heatid="20005">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:04.16" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="128" birthdate="2014-01-01" gender="M" lastname="Michalke" firstname="Max-Leon" license="0">
              <RESULTS>
                <RESULT resultid="351" eventid="8" swimtime="00:01:25.32" lane="4" heatid="8001" />
                <RESULT resultid="352" eventid="15" swimtime="00:00:38.31" lane="7" heatid="15002" />
                <RESULT resultid="353" eventid="21" swimtime="00:03:09.79" lane="2" heatid="21001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:35.62" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="129" birthdate="2013-01-01" gender="M" lastname="Hartmann" firstname="Paul" license="0">
              <RESULTS>
                <RESULT resultid="354" eventid="8" swimtime="00:01:14.98" reactiontime="+94" lane="7" heatid="8003" />
                <RESULT resultid="355" eventid="15" swimtime="00:00:35.56" lane="4" heatid="15003" />
                <RESULT resultid="356" eventid="21" swimtime="00:02:48.16" lane="5" heatid="21001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:21.31" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="130" birthdate="1964-01-01" gender="F" lastname="Saliger" firstname="Petra" license="0">
              <RESULTS>
                <RESULT resultid="357" eventid="7" swimtime="00:01:15.43" reactiontime="+88" lane="6" heatid="7004" />
                <RESULT resultid="358" eventid="14" swimtime="00:00:34.49" lane="3" heatid="14004" />
                <RESULT resultid="359" eventid="18" swimtime="00:01:33.03" lane="3" heatid="18001" />
                <RESULT resultid="360" eventid="22" swimtime="00:07:24.44" lane="8" heatid="22001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:39.59" />
                    <SPLIT distance="200" swimtime="00:03:34.63" />
                    <SPLIT distance="300" swimtime="00:05:31.25" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="131" birthdate="1953-01-01" gender="F" lastname="Reuter" firstname="Renate" license="0">
              <RESULTS>
                <RESULT resultid="361" eventid="7" status="DNS" swimtime="00:00:00.00" lane="8" heatid="7002" />
                <RESULT resultid="362" eventid="14" swimtime="00:00:42.46" lane="1" heatid="14002" />
                <RESULT resultid="363" eventid="18" status="DNS" swimtime="00:00:00.00" lane="6" heatid="18001" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="132" birthdate="1959-01-01" gender="M" lastname="Senf" firstname="Rüdiger" license="0">
              <RESULTS>
                <RESULT resultid="364" eventid="2" swimtime="00:05:14.60" reactiontime="+99" lane="4" heatid="2002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:14.24" />
                    <SPLIT distance="200" swimtime="00:02:35.99" />
                    <SPLIT distance="300" swimtime="00:03:57.99" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="365" eventid="8" swimtime="00:01:05.47" lane="2" heatid="8005" />
                <RESULT resultid="366" eventid="12" swimtime="00:00:30.14" lane="5" heatid="12001" />
                <RESULT resultid="367" eventid="15" swimtime="00:00:30.36" lane="3" heatid="15005" />
                <RESULT resultid="368" eventid="21" swimtime="00:02:34.82" lane="4" heatid="21003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:13.15" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="133" birthdate="2008-01-01" gender="F" lastname="Steinert" firstname="Sara-Marie" license="0">
              <RESULTS>
                <RESULT resultid="369" eventid="7" swimtime="00:01:53.47" lane="4" heatid="7001" />
                <RESULT resultid="370" eventid="14" swimtime="00:00:41.34" lane="5" heatid="14001" />
                <RESULT resultid="371" eventid="20" swimtime="00:03:35.04" lane="1" heatid="20002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:38.87" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="134" birthdate="1972-01-01" gender="M" lastname="Gräf" firstname="Sven" license="0">
              <RESULTS>
                <RESULT resultid="372" eventid="12" swimtime="00:00:23.27" lane="4" heatid="12002" />
                <RESULT resultid="373" eventid="15" swimtime="00:00:20.28" lane="8" heatid="15009" />
                <RESULT resultid="374" eventid="19" swimtime="00:00:42.86" lane="3" heatid="19002" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="135" birthdate="2010-01-01" gender="F" lastname="Martin" firstname="Theresa" license="0">
              <RESULTS>
                <RESULT resultid="375" eventid="1" swimtime="00:05:18.85" reactiontime="+94" lane="6" heatid="1002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:12.62" />
                    <SPLIT distance="200" swimtime="00:02:36.06" />
                    <SPLIT distance="300" swimtime="00:04:01.75" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="376" eventid="7" swimtime="00:01:04.78" reactiontime="+97" lane="6" heatid="7005" />
                <RESULT resultid="377" eventid="14" swimtime="00:00:29.08" lane="5" heatid="14005" />
                <RESULT resultid="378" eventid="20" swimtime="00:02:27.35" lane="4" heatid="20004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:10.02" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="136" birthdate="2012-01-01" gender="F" lastname="Riedel" firstname="Valentina" license="0">
              <RESULTS>
                <RESULT resultid="379" eventid="7" swimtime="00:01:20.21" lane="3" heatid="7002" />
                <RESULT resultid="380" eventid="14" swimtime="00:00:35.30" lane="7" heatid="14003" />
                <RESULT resultid="381" eventid="20" swimtime="00:03:04.57" reactiontime="+60" lane="3" heatid="20002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:31.73" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="137" birthdate="2013-01-01" gender="M" lastname="Kad" firstname="Vincent" license="0">
              <RESULTS>
                <RESULT resultid="382" eventid="8" swimtime="00:01:26.89" lane="1" heatid="8002" />
                <RESULT resultid="383" eventid="15" swimtime="00:00:39.17" lane="5" heatid="15002" />
                <RESULT resultid="384" eventid="21" swimtime="00:03:20.52" lane="3" heatid="21001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:40.91" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY number="1" gender="X" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="321" eventid="13" swimtime="00:02:01.64" lane="1" heatid="13002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:02.54" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="128" number="1" />
                    <RELAYPOSITION athleteid="127" number="2" />
                    <RELAYPOSITION athleteid="129" number="3" />
                    <RELAYPOSITION athleteid="123" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="2" gender="F" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="322" eventid="24" swimtime="00:04:12.70" lane="7" heatid="24002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:58.71" />
                    <SPLIT distance="200" swimtime="00:02:05.43" />
                    <SPLIT distance="300" swimtime="00:03:23.59" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="135" number="1" />
                    <RELAYPOSITION athleteid="127" number="2" />
                    <RELAYPOSITION athleteid="125" number="3" />
                    <RELAYPOSITION athleteid="123" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="3" gender="X" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="323" eventid="13" swimtime="00:02:17.63" lane="4" heatid="13001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:05.44" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="132" number="1" />
                    <RELAYPOSITION athleteid="130" number="2" />
                    <RELAYPOSITION athleteid="131" number="3" />
                    <RELAYPOSITION athleteid="121" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB name="Tauchsport Döbeln" nation="GER" region="20" code="154104000">
          <ATHLETES>
            <ATHLETE athleteid="10" birthdate="2006-01-01" gender="M" lastname="Noack" firstname="Christopher" license="0">
              <RESULTS>
                <RESULT resultid="39" eventid="6" status="DSQ" swimtime="00:00:26.84" lane="4" heatid="6001" comment="Gesicht aus dem Wasser bei 30 Meter." />
                <RESULT resultid="40" eventid="8" swimtime="00:00:55.46" lane="2" heatid="8006" />
                <RESULT resultid="41" eventid="15" swimtime="00:00:24.14" lane="4" heatid="15006" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="11" birthdate="1973-01-01" gender="M" lastname="Winkler" firstname="Daniel" license="0">
              <RESULTS>
                <RESULT resultid="42" eventid="6" swimtime="00:00:21.36" lane="1" heatid="6003" />
                <RESULT resultid="43" eventid="8" swimtime="00:00:52.31" lane="8" heatid="8007" />
                <RESULT resultid="44" eventid="12" status="DSQ" swimtime="00:00:25.42" lane="2" heatid="12002" comment="Falscher Start." />
                <RESULT resultid="45" eventid="15" swimtime="00:00:23.56" lane="3" heatid="15007" />
                <RESULT resultid="46" eventid="19" swimtime="00:00:51.22" lane="4" heatid="19001" />
                <RESULT resultid="47" eventid="21" swimtime="00:02:05.70" lane="7" heatid="21005">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:59.03" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="12" birthdate="2003-01-01" gender="M" lastname="Elenkow" firstname="Felix" license="0">
              <RESULTS>
                <RESULT resultid="48" eventid="6" swimtime="00:00:18.80" lane="1" heatid="6004" />
                <RESULT resultid="49" eventid="8" swimtime="00:00:45.99" reactiontime="+93" lane="8" heatid="8008" />
                <RESULT resultid="50" eventid="15" swimtime="00:00:20.72" lane="2" heatid="15008" />
                <RESULT resultid="51" eventid="19" swimtime="00:00:46.39" lane="2" heatid="19002" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="13" birthdate="1962-01-01" gender="M" lastname="Muth" firstname="Henrik" license="0">
              <RESULTS>
                <RESULT resultid="52" eventid="2" swimtime="00:04:53.96" lane="7" heatid="2003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:06.46" />
                    <SPLIT distance="200" swimtime="00:02:22.37" />
                    <SPLIT distance="300" swimtime="00:03:39.08" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="53" eventid="6" swimtime="00:00:20.74" lane="2" heatid="6003" />
                <RESULT resultid="54" eventid="8" swimtime="00:00:51.84" lane="4" heatid="8006" />
                <RESULT resultid="55" eventid="10" swimtime="00:10:13.44" lane="1" heatid="10001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:09.36" />
                    <SPLIT distance="200" swimtime="00:02:26.15" />
                    <SPLIT distance="300" swimtime="00:03:45.13" />
                    <SPLIT distance="400" swimtime="00:05:03.71" />
                    <SPLIT distance="500" swimtime="00:06:23.16" />
                    <SPLIT distance="600" swimtime="00:07:43.22" />
                    <SPLIT distance="700" swimtime="00:09:02.14" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="56" eventid="15" swimtime="00:00:25.07" lane="5" heatid="15006" />
                <RESULT resultid="57" eventid="19" swimtime="00:00:49.16" lane="8" heatid="19002" />
                <RESULT resultid="58" eventid="21" swimtime="00:02:09.78" lane="4" heatid="21004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:02.20" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="59" eventid="23" swimtime="00:04:34.56" lane="1" heatid="23001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:01.17" />
                    <SPLIT distance="200" swimtime="00:02:12.46" />
                    <SPLIT distance="300" swimtime="00:03:24.75" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="14" birthdate="2006-01-01" gender="F" lastname="Elenkow" firstname="Johanna" license="0">
              <RESULTS>
                <RESULT resultid="60" eventid="5" swimtime="00:00:30.35" lane="6" heatid="5001" />
                <RESULT resultid="61" eventid="7" swimtime="00:01:03.28" lane="5" heatid="7005" />
                <RESULT resultid="62" eventid="14" swimtime="00:00:28.77" lane="3" heatid="14006" />
                <RESULT resultid="63" eventid="20" swimtime="00:02:30.49" lane="3" heatid="20003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:08.22" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="15" birthdate="1972-01-01" gender="M" lastname="Schuricht" firstname="Oliver" license="0">
              <RESULTS>
                <RESULT resultid="64" eventid="12" swimtime="00:00:24.90" lane="7" heatid="12002" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="Tauchsportclub Erfurt e.V." nation="GER" region="35" code="0">
          <ATHLETES>
            <ATHLETE athleteid="66" birthdate="2010-01-01" gender="F" lastname="Abe" firstname="Adina" license="0">
              <RESULTS>
                <RESULT resultid="660" eventid="3" swimtime="00:00:23.31" lane="4" heatid="3001" />
                <RESULT resultid="661" eventid="7" swimtime="00:00:51.35" lane="7" heatid="7008" />
                <RESULT resultid="662" eventid="14" swimtime="00:00:23.56" lane="8" heatid="14009" />
                <RESULT resultid="663" eventid="20" swimtime="00:01:55.45" lane="1" heatid="20006">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:56.06" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="67" birthdate="2009-01-01" gender="F" lastname="Zitzmann" firstname="Annalena" license="0">
              <RESULTS>
                <RESULT resultid="664" eventid="5" swimtime="00:00:22.79" lane="6" heatid="5002" />
                <RESULT resultid="665" eventid="7" swimtime="00:00:51.88" reactiontime="+93" lane="5" heatid="7007" />
                <RESULT resultid="666" eventid="14" swimtime="00:00:23.46" lane="6" heatid="14009" />
                <RESULT resultid="667" eventid="18" swimtime="00:00:54.53" lane="1" heatid="18003" />
                <RESULT resultid="668" eventid="20" swimtime="00:02:01.23" reactiontime="+98" lane="3" heatid="20005">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:57.86" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="68" birthdate="2011-01-01" gender="F" lastname="Behrmann" firstname="Fine Erna" license="0">
              <RESULTS>
                <RESULT resultid="669" eventid="3" swimtime="00:00:30.41" lane="6" heatid="3001" />
                <RESULT resultid="670" eventid="7" swimtime="00:01:03.84" lane="4" heatid="7005" />
                <RESULT resultid="671" eventid="14" swimtime="00:00:28.77" lane="8" heatid="14007" />
                <RESULT resultid="672" eventid="20" swimtime="00:02:20.04" lane="7" heatid="20004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:06.42" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="69" birthdate="2009-01-01" gender="M" lastname="Artschwager" firstname="Gustaf" license="0">
              <RESULTS>
                <RESULT resultid="673" eventid="2" swimtime="00:04:56.71" lane="2" heatid="2003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:06.40" />
                    <SPLIT distance="200" swimtime="00:02:23.50" />
                    <SPLIT distance="300" swimtime="00:03:41.88" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="674" eventid="8" swimtime="00:01:04.02" lane="5" heatid="8005" />
                <RESULT resultid="675" eventid="15" swimtime="00:00:29.81" lane="7" heatid="15006" />
                <RESULT resultid="676" eventid="21" swimtime="00:02:13.97" reactiontime="+95" lane="5" heatid="21004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:04.55" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="71" birthdate="2010-01-01" gender="M" lastname="Schmidt" firstname="Jakob" license="0">
              <RESULTS>
                <RESULT resultid="677" eventid="2" swimtime="00:06:17.35" reactiontime="+91" lane="5" heatid="2001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:20.33" />
                    <SPLIT distance="200" swimtime="00:02:59.65" />
                    <SPLIT distance="300" swimtime="00:04:41.46" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="678" eventid="8" swimtime="00:01:24.98" reactiontime="+89" lane="5" heatid="8003" />
                <RESULT resultid="679" eventid="15" swimtime="00:00:36.08" lane="3" heatid="15004" />
                <RESULT resultid="680" eventid="21" swimtime="00:02:56.45" reactiontime="+85" lane="5" heatid="21002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:24.90" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="72" birthdate="2010-01-01" gender="M" lastname="Hochstein" firstname="Jean Paul" license="0">
              <RESULTS>
                <RESULT resultid="681" eventid="4" swimtime="00:00:29.13" lane="5" heatid="4001" />
                <RESULT resultid="682" eventid="8" swimtime="00:00:58.89" reactiontime="+85" lane="4" heatid="8005" />
                <RESULT resultid="683" eventid="15" swimtime="00:00:26.15" lane="3" heatid="15006" />
                <RESULT resultid="684" eventid="21" swimtime="00:02:16.12" reactiontime="+95" lane="7" heatid="21004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:06.70" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="73" birthdate="2006-01-01" gender="M" lastname="Leipold" firstname="Marek" license="0">
              <RESULTS>
                <RESULT resultid="689" eventid="6" swimtime="00:00:15.54" lane="4" heatid="6004" />
                <RESULT resultid="690" eventid="8" swimtime="00:00:37.22" reactiontime="+88" lane="4" heatid="8008" />
                <RESULT resultid="691" eventid="15" swimtime="00:00:16.51" lane="4" heatid="15009" />
                <RESULT resultid="692" eventid="21" swimtime="00:01:28.00" reactiontime="+90" lane="4" heatid="21006">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:40.38" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="74" birthdate="2009-01-01" gender="F" lastname="Blumenstein" firstname="Martha" license="0">
              <RESULTS>
                <RESULT resultid="693" eventid="1" swimtime="00:04:29.98" reactiontime="+91" lane="3" heatid="1003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:01.61" />
                    <SPLIT distance="200" swimtime="00:02:12.30" />
                    <SPLIT distance="300" swimtime="00:03:23.30" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="694" eventid="7" swimtime="00:00:54.44" reactiontime="+89" lane="5" heatid="7006" />
                <RESULT resultid="695" eventid="14" swimtime="00:00:23.98" lane="6" heatid="14008" />
                <RESULT resultid="696" eventid="20" swimtime="00:02:06.29" lane="2" heatid="20005">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:01.19" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="75" birthdate="1979-01-01" gender="F" lastname="Leipold" firstname="Steffi" license="0">
              <RESULTS>
                <RESULT resultid="697" eventid="5" swimtime="00:00:25.03" lane="5" heatid="5001" />
                <RESULT resultid="698" eventid="14" swimtime="00:00:25.89" lane="4" heatid="14007" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="76" birthdate="1963-01-01" gender="F" lastname="Tiszold" firstname="Ursula" license="0">
              <RESULTS>
                <RESULT resultid="699" eventid="1" swimtime="00:05:43.41" lane="3" heatid="1002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:14.18" />
                    <SPLIT distance="200" swimtime="00:02:42.07" />
                    <SPLIT distance="300" swimtime="00:04:14.96" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="700" eventid="5" swimtime="00:00:38.18" lane="1" heatid="5001" />
                <RESULT resultid="701" eventid="7" swimtime="00:01:09.76" lane="2" heatid="7005" />
                <RESULT resultid="702" eventid="11" swimtime="00:00:31.94" lane="7" heatid="11001" />
                <RESULT resultid="703" eventid="14" swimtime="00:00:31.82" lane="4" heatid="14005" />
                <RESULT resultid="704" eventid="20" swimtime="00:02:43.57" lane="1" heatid="20004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:14.72" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="293" birthdate="2006-01-01" gender="F" lastname="Heinitz" firstname="Leonor" license="0">
              <RESULTS>
                <RESULT resultid="685" eventid="5" swimtime="00:00:22.14" lane="5" heatid="5002" />
                <RESULT resultid="686" eventid="7" swimtime="00:00:53.58" lane="3" heatid="7007" />
                <RESULT resultid="687" eventid="14" swimtime="00:00:23.85" lane="3" heatid="14008" />
                <RESULT resultid="688" eventid="18" swimtime="00:00:52.59" lane="5" heatid="18002" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY number="1" gender="X" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="" />
            <RELAY number="2" gender="F" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="659" eventid="24" swimtime="00:03:44.78" lane="2" heatid="24002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:53.19" />
                    <SPLIT distance="200" swimtime="00:01:51.14" />
                    <SPLIT distance="300" swimtime="00:02:52.99" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="67" number="1" />
                    <RELAYPOSITION athleteid="74" number="2" />
                    <RELAYPOSITION athleteid="68" number="3" />
                    <RELAYPOSITION athleteid="66" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" gender="X" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="658" eventid="13" swimtime="00:01:42.06" lane="7" heatid="13002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:49.50" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="72" number="1" />
                    <RELAYPOSITION athleteid="67" number="2" />
                    <RELAYPOSITION athleteid="69" number="3" />
                    <RELAYPOSITION athleteid="66" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB name="TC Chemie Greiz e.V." nation="GER" region="35" code="174117">
          <ATHLETES>
            <ATHLETE athleteid="33" birthdate="2006-01-01" gender="F" lastname="Frauenfelder" firstname="Anneliese" license="0">
              <RESULTS>
                <RESULT resultid="86" eventid="5" swimtime="00:00:21.61" lane="6" heatid="5003" />
                <RESULT resultid="87" eventid="7" swimtime="00:00:50.10" reactiontime="+94" lane="4" heatid="7008" />
                <RESULT resultid="88" eventid="14" swimtime="00:00:23.24" lane="3" heatid="14009" />
                <RESULT resultid="89" eventid="18" swimtime="00:00:48.86" lane="8" heatid="18004" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="35" birthdate="2011-01-01" gender="F" lastname="Volger" firstname="Eva" license="0">
              <RESULTS>
                <RESULT resultid="93" eventid="1" swimtime="00:05:59.08" reactiontime="+99" lane="7" heatid="1002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:21.62" />
                    <SPLIT distance="200" swimtime="00:02:53.86" />
                    <SPLIT distance="300" swimtime="00:04:28.86" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="94" eventid="7" swimtime="00:01:14.86" reactiontime="+90" lane="4" heatid="7003" />
                <RESULT resultid="95" eventid="14" swimtime="00:00:33.35" lane="2" heatid="14004" />
                <RESULT resultid="96" eventid="20" swimtime="00:02:47.31" reactiontime="+97" lane="1" heatid="20003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:20.37" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="36" birthdate="2016-01-01" gender="F" lastname="Volger" firstname="Lea" license="0">
              <RESULTS>
                <RESULT resultid="97" eventid="7" swimtime="00:01:25.33" lane="1" heatid="7002" />
                <RESULT resultid="98" eventid="14" swimtime="00:00:39.11" lane="2" heatid="14002" />
                <RESULT resultid="99" eventid="20" swimtime="00:03:24.89" lane="6" heatid="20002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:45.55" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="37" birthdate="2013-01-01" gender="F" lastname="Jutzenka" firstname="Leonie" license="0">
              <RESULTS>
                <RESULT resultid="100" eventid="1" swimtime="00:06:46.51" lane="1" heatid="1002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:36.09" />
                    <SPLIT distance="200" swimtime="00:03:21.09" />
                    <SPLIT distance="300" swimtime="00:05:07.20" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="101" eventid="7" swimtime="00:01:27.57" lane="5" heatid="7002" />
                <RESULT resultid="102" eventid="14" swimtime="00:00:37.82" lane="3" heatid="14002" />
                <RESULT resultid="103" eventid="20" swimtime="00:01:30.05" lane="4" heatid="20005">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:03:09.07" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="38" birthdate="2014-01-01" gender="F" lastname="Blei" firstname="Lina" license="0">
              <RESULTS>
                <RESULT resultid="104" eventid="7" status="DNS" swimtime="00:00:00.00" lane="3" heatid="7001" />
                <RESULT resultid="105" eventid="14" status="DNS" swimtime="00:00:00.00" lane="4" heatid="14001" />
                <RESULT resultid="106" eventid="20" status="DNS" swimtime="00:00:00.00" lane="4" heatid="20001" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="39" birthdate="2008-01-01" gender="M" lastname="Berger" firstname="Louis" license="0">
              <RESULTS>
                <RESULT resultid="107" eventid="2" status="DNS" swimtime="00:00:00.00" lane="6" heatid="2004" />
                <RESULT resultid="108" eventid="15" status="DNS" swimtime="00:00:00.00" lane="5" heatid="15008" />
                <RESULT resultid="109" eventid="21" status="DNS" swimtime="00:00:00.00" lane="2" heatid="21006" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="40" birthdate="2005-01-01" gender="F" lastname="Kupka" firstname="Miriam" license="0">
              <RESULTS>
                <RESULT resultid="110" eventid="1" swimtime="00:03:58.20" reactiontime="+93" lane="1" heatid="1005">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:55.28" />
                    <SPLIT distance="200" swimtime="00:01:56.87" />
                    <SPLIT distance="300" swimtime="00:02:59.03" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="111" eventid="7" swimtime="00:00:46.78" reactiontime="+91" lane="5" heatid="7009" />
                <RESULT resultid="112" eventid="14" swimtime="00:00:20.93" lane="8" heatid="14011" />
                <RESULT resultid="113" eventid="20" swimtime="00:01:50.44" reactiontime="+96" lane="4" heatid="20006">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:53.27" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="41" birthdate="2015-01-01" gender="M" lastname="Kießling" firstname="Moritz" license="0">
              <RESULTS>
                <RESULT resultid="114" eventid="8" swimtime="00:02:03.86" reactiontime="+99" lane="3" heatid="8001" />
                <RESULT resultid="115" eventid="15" status="DSQ" swimtime="00:00:40.60" lane="4" heatid="15001" comment="Falscher Start." />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="42" birthdate="1974-01-01" gender="M" lastname="Kühn" firstname="Ronald" license="0">
              <RESULTS>
                <RESULT resultid="116" eventid="6" swimtime="00:00:21.42" lane="3" heatid="6003" />
                <RESULT resultid="117" eventid="8" swimtime="00:00:56.34" lane="1" heatid="8007" />
                <RESULT resultid="118" eventid="15" swimtime="00:00:25.12" lane="7" heatid="15007" />
                <RESULT resultid="119" eventid="21" swimtime="00:02:10.98" reactiontime="+95" lane="1" heatid="21005">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:02.38" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="43" birthdate="2011-01-01" gender="F" lastname="Leonhardt" firstname="Ronja" license="0">
              <RESULTS>
                <RESULT resultid="120" eventid="1" status="DNS" swimtime="00:00:00.00" lane="2" heatid="1002" />
                <RESULT resultid="121" eventid="9" status="DNS" swimtime="00:00:00.00" lane="3" heatid="9001" />
                <RESULT resultid="122" eventid="14" status="DNS" swimtime="00:00:00.00" lane="5" heatid="14004" />
                <RESULT resultid="123" eventid="20" status="DNS" swimtime="00:00:00.00" lane="4" heatid="20003" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="44" birthdate="2013-01-01" gender="M" lastname="Robenz" firstname="Ronny Jason" license="0">
              <RESULTS>
                <RESULT resultid="124" eventid="2" swimtime="00:05:45.52" lane="2" heatid="2002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:19.11" />
                    <SPLIT distance="200" swimtime="00:02:50.16" />
                    <SPLIT distance="300" swimtime="00:04:19.52" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="125" eventid="8" swimtime="00:01:15.85" reactiontime="+94" lane="7" heatid="8004" />
                <RESULT resultid="126" eventid="15" swimtime="00:00:33.28" lane="1" heatid="15004" />
                <RESULT resultid="127" eventid="21" swimtime="00:02:40.23" reactiontime="+98" lane="4" heatid="21002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:17.88" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="45" birthdate="2011-01-01" gender="F" lastname="Klar" firstname="Sophia" license="0">
              <RESULTS>
                <RESULT resultid="128" eventid="3" swimtime="00:00:32.13" lane="2" heatid="3001" />
                <RESULT resultid="129" eventid="9" swimtime="00:14:08.91" lane="5" heatid="9001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:32.39" />
                    <SPLIT distance="200" swimtime="00:03:21.39" />
                    <SPLIT distance="300" swimtime="00:05:09.83" />
                    <SPLIT distance="400" swimtime="00:07:01.06" />
                    <SPLIT distance="500" swimtime="00:08:51.54" />
                    <SPLIT distance="600" swimtime="00:10:45.56" />
                    <SPLIT distance="700" swimtime="00:12:32.15" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="130" eventid="14" swimtime="00:00:31.17" lane="6" heatid="14005" />
                <RESULT resultid="131" eventid="18" swimtime="00:01:21.04" lane="5" heatid="18001" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="46" birthdate="2016-01-01" gender="M" lastname="Hierold" firstname="Theodor" license="0">
              <RESULTS>
                <RESULT resultid="132" eventid="8" swimtime="00:01:34.00" lane="8" heatid="8002" />
                <RESULT resultid="133" eventid="15" swimtime="00:00:39.74" lane="4" heatid="15002" />
                <RESULT resultid="134" eventid="21" swimtime="00:03:29.04" lane="4" heatid="21001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:41.41" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="47" birthdate="2000-01-01" gender="M" lastname="Kupka" firstname="Titus" license="0">
              <RESULTS>
                <RESULT resultid="135" eventid="6" swimtime="00:00:17.53" lane="3" heatid="6004" />
                <RESULT resultid="136" eventid="8" swimtime="00:00:43.40" reactiontime="+91" lane="2" heatid="8008" />
                <RESULT resultid="137" eventid="15" swimtime="00:00:19.27" lane="4" heatid="15008" />
                <RESULT resultid="138" eventid="19" swimtime="00:00:42.54" lane="4" heatid="19002" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="48" birthdate="2014-01-01" gender="M" lastname="Volger" firstname="Tom" license="0">
              <RESULTS>
                <RESULT resultid="139" eventid="2" swimtime="00:06:02.95" reactiontime="+98" lane="4" heatid="2001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:21.29" />
                    <SPLIT distance="200" swimtime="00:02:53.36" />
                    <SPLIT distance="300" swimtime="00:04:28.90" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="140" eventid="8" swimtime="00:01:19.41" reactiontime="+97" lane="6" heatid="8003" />
                <RESULT resultid="141" eventid="15" swimtime="00:00:34.56" lane="2" heatid="15003" />
                <RESULT resultid="142" eventid="21" swimtime="00:02:46.68" reactiontime="+92" lane="6" heatid="21002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:21.08" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="49" birthdate="2012-01-01" gender="M" lastname="Sochynskyi" firstname="Vadym" license="0">
              <RESULTS>
                <RESULT resultid="143" eventid="2" swimtime="00:05:28.48" reactiontime="+94" lane="6" heatid="2002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:16.76" />
                    <SPLIT distance="200" swimtime="00:02:42.65" />
                    <SPLIT distance="300" swimtime="00:04:07.54" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="144" eventid="8" swimtime="00:01:07.67" reactiontime="+87" lane="2" heatid="8004" />
                <RESULT resultid="145" eventid="15" swimtime="00:00:30.47" lane="1" heatid="15005" />
                <RESULT resultid="146" eventid="21" swimtime="00:02:33.43" reactiontime="+91" lane="1" heatid="21003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:16.44" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="TC Delitzsch" nation="GER" region="20" code="0">
          <ATHLETES>
            <ATHLETE athleteid="148" birthdate="1999-01-01" gender="F" lastname="Gusmanov" firstname="Jil" license="0">
              <RESULTS>
                <RESULT resultid="413" eventid="1" swimtime="00:04:46.67" lane="7" heatid="1003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:07.19" />
                    <SPLIT distance="200" swimtime="00:02:19.11" />
                    <SPLIT distance="300" swimtime="00:03:33.04" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="414" eventid="9" swimtime="00:09:56.65" lane="4" heatid="9001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:10.42" />
                    <SPLIT distance="200" swimtime="00:02:24.71" />
                    <SPLIT distance="300" swimtime="00:03:40.12" />
                    <SPLIT distance="400" swimtime="00:04:55.29" />
                    <SPLIT distance="500" swimtime="00:06:10.88" />
                    <SPLIT distance="600" swimtime="00:07:27.37" />
                    <SPLIT distance="700" swimtime="00:08:41.85" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="415" eventid="20" swimtime="00:02:17.43" lane="6" heatid="20004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:05.17" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="149" birthdate="2011-01-01" gender="F" lastname="Schönherr" firstname="Nina" license="0">
              <RESULTS>
                <RESULT resultid="416" eventid="3" swimtime="00:00:27.12" lane="1" heatid="3001" />
                <RESULT resultid="417" eventid="7" swimtime="00:00:57.48" reactiontime="+94" lane="6" heatid="7006" />
                <RESULT resultid="418" eventid="14" swimtime="00:00:26.97" lane="5" heatid="14007" />
                <RESULT resultid="419" eventid="18" swimtime="00:01:01.68" lane="4" heatid="18001" />
                <RESULT resultid="420" eventid="20" swimtime="00:02:17.20" reactiontime="+80" lane="3" heatid="20004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:06.68" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="150" birthdate="2011-01-01" gender="M" lastname="Becker" firstname="Pepe Milan" license="0">
              <RESULTS>
                <RESULT resultid="421" eventid="4" swimtime="00:00:30.63" lane="3" heatid="4001" />
                <RESULT resultid="422" eventid="8" swimtime="00:01:00.52" reactiontime="+95" lane="1" heatid="8004" />
                <RESULT resultid="423" eventid="15" swimtime="00:00:26.38" lane="4" heatid="15005" />
                <RESULT resultid="424" eventid="19" swimtime="00:01:10.16" lane="7" heatid="19001" />
                <RESULT resultid="425" eventid="21" swimtime="00:02:16.51" reactiontime="+94" lane="3" heatid="21003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:05.67" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="TC fez Berlin" nation="GER" region="21" code="34113000">
          <ATHLETES>
            <ATHLETE athleteid="195" birthdate="2006-01-01" gender="M" lastname="Schlobohm" firstname="Enrico" license="3411">
              <RESULTS>
                <RESULT resultid="535" eventid="6" swimtime="00:00:17.41" lane="2" heatid="6004" />
                <RESULT resultid="536" eventid="8" swimtime="00:00:45.02" reactiontime="+84" lane="7" heatid="8008" />
                <RESULT resultid="537" eventid="15" swimtime="00:00:19.83" lane="3" heatid="15008" />
                <RESULT resultid="538" eventid="21" swimtime="00:01:46.68" lane="7" heatid="21006">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:49.59" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="196" birthdate="1996-01-01" gender="M" lastname="Schustek" firstname="Fabian" license="0">
              <RESULTS>
                <RESULT resultid="539" eventid="6" swimtime="00:00:17.77" lane="7" heatid="6004" />
                <RESULT resultid="540" eventid="8" swimtime="00:00:41.81" reactiontime="+89" lane="6" heatid="8008" />
                <RESULT resultid="651" eventid="15" swimtime="00:00:19.11" lane="7" heatid="15009" />
                <RESULT resultid="541" eventid="19" swimtime="00:00:42.99" lane="6" heatid="19002" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="197" birthdate="2002-01-01" gender="F" lastname="Schikora" firstname="Johanna" license="0">
              <RESULTS>
                <RESULT resultid="543" eventid="1" swimtime="00:03:23.30" reactiontime="+99" lane="4" heatid="1005">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:49.65" />
                    <SPLIT distance="200" swimtime="00:01:40.85" />
                    <SPLIT distance="300" swimtime="00:02:32.76" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="544" eventid="7" swimtime="00:00:44.49" reactiontime="+97" lane="6" heatid="7010" />
                <RESULT resultid="545" eventid="14" swimtime="00:00:21.25" lane="5" heatid="14010" />
                <RESULT resultid="546" eventid="20" swimtime="00:01:34.53" reactiontime="+98" lane="4" heatid="20007">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:46.57" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="198" birthdate="2006-01-01" gender="F" lastname="Zobel" firstname="Juliane" license="341100319">
              <RESULTS>
                <RESULT resultid="547" eventid="1" status="DSQ" swimtime="00:04:02.25" reactiontime="+88" lane="5" heatid="1004" comment="Tauchzüge bei ca. 200 Meter.">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:55.14" />
                    <SPLIT distance="200" swimtime="00:01:56.91" />
                    <SPLIT distance="300" swimtime="00:03:00.70" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="548" eventid="5" swimtime="00:00:21.71" lane="4" heatid="5002" />
                <RESULT resultid="549" eventid="7" swimtime="00:00:49.74" reactiontime="+86" lane="5" heatid="7008" />
                <RESULT resultid="550" eventid="14" swimtime="00:00:21.90" lane="8" heatid="14010" />
                <RESULT resultid="551" eventid="18" swimtime="00:00:49.41" lane="7" heatid="18003" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="199" birthdate="2005-01-01" gender="F" lastname="Gawenda" firstname="Lara" license="0">
              <RESULTS>
                <RESULT resultid="552" eventid="5" status="DNS" swimtime="00:00:00.00" lane="5" heatid="5004" />
                <RESULT resultid="553" eventid="7" status="DNS" swimtime="00:00:00.00" lane="5" heatid="7010" />
                <RESULT resultid="554" eventid="14" status="DNS" swimtime="00:00:00.00" lane="5" heatid="14011" />
                <RESULT resultid="555" eventid="20" status="DNS" swimtime="00:00:00.00" lane="5" heatid="20007" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="200" birthdate="2008-01-01" gender="F" lastname="Sunagatova" firstname="Milana" license="0">
              <RESULTS>
                <RESULT resultid="556" eventid="1" swimtime="00:03:47.28" lane="7" heatid="1005">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:52.80" />
                    <SPLIT distance="200" swimtime="00:01:51.04" />
                    <SPLIT distance="300" swimtime="00:02:49.49" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="557" eventid="7" swimtime="00:00:47.61" lane="6" heatid="7009" />
                <RESULT resultid="558" eventid="9" swimtime="00:08:05.55" lane="3" heatid="9002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:55.41" />
                    <SPLIT distance="200" swimtime="00:01:56.50" />
                    <SPLIT distance="300" swimtime="00:02:58.66" />
                    <SPLIT distance="400" swimtime="00:04:00.97" />
                    <SPLIT distance="500" swimtime="00:05:02.62" />
                    <SPLIT distance="600" swimtime="00:06:04.21" />
                    <SPLIT distance="700" swimtime="00:07:06.37" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="559" eventid="14" swimtime="00:00:22.05" lane="5" heatid="14009" />
                <RESULT resultid="560" eventid="20" swimtime="00:01:45.38" lane="5" heatid="20006">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:50.98" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="201" birthdate="2006-01-01" gender="F" lastname="Ahnert" firstname="Paula" license="0">
              <RESULTS>
                <RESULT resultid="561" eventid="1" swimtime="00:03:57.42" reactiontime="+88" lane="6" heatid="1005">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:53.92" />
                    <SPLIT distance="200" swimtime="00:01:53.01" />
                    <SPLIT distance="300" swimtime="00:02:54.65" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="562" eventid="5" swimtime="00:00:19.80" lane="4" heatid="5003" />
                <RESULT resultid="563" eventid="7" swimtime="00:00:46.31" reactiontime="+87" lane="1" heatid="7010" />
                <RESULT resultid="564" eventid="9" swimtime="00:08:00.51" reactiontime="+85" lane="4" heatid="9002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:55.30" />
                    <SPLIT distance="200" swimtime="00:01:55.52" />
                    <SPLIT distance="300" swimtime="00:02:56.22" />
                    <SPLIT distance="400" swimtime="00:03:57.97" />
                    <SPLIT distance="500" swimtime="00:04:58.76" />
                    <SPLIT distance="600" swimtime="00:06:00.06" />
                    <SPLIT distance="700" swimtime="00:07:00.76" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="565" eventid="14" swimtime="00:00:21.07" lane="3" heatid="14010" />
                <RESULT resultid="566" eventid="20" swimtime="00:01:47.63" reactiontime="+91" lane="1" heatid="20007">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:50.35" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="202" birthdate="2002-01-01" gender="M" lastname="Lebeau" firstname="Remy" license="0">
              <RESULTS>
                <RESULT resultid="567" eventid="2" swimtime="00:03:21.75" reactiontime="+95" lane="5" heatid="2004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:47.34" />
                    <SPLIT distance="200" swimtime="00:01:38.83" />
                    <SPLIT distance="300" swimtime="00:02:31.07" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="568" eventid="8" swimtime="00:00:43.47" reactiontime="+97" lane="3" heatid="8008" />
                <RESULT resultid="569" eventid="15" swimtime="00:00:19.66" lane="1" heatid="15009" />
                <RESULT resultid="570" eventid="21" swimtime="00:01:33.90" reactiontime="+96" lane="5" heatid="21006">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:45.00" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="203" birthdate="2006-01-01" gender="M" lastname="Patge" firstname="Rufus" license="3411">
              <RESULTS>
                <RESULT resultid="571" eventid="2" swimtime="00:04:01.29" reactiontime="+91" lane="2" heatid="2004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:52.58" />
                    <SPLIT distance="200" swimtime="00:01:52.32" />
                    <SPLIT distance="300" swimtime="00:02:53.96" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="572" eventid="10" swimtime="00:08:24.88" reactiontime="+95" lane="6" heatid="10001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:55.32" />
                    <SPLIT distance="200" swimtime="00:01:58.87" />
                    <SPLIT distance="300" swimtime="00:03:03.77" />
                    <SPLIT distance="400" swimtime="00:04:09.66" />
                    <SPLIT distance="500" swimtime="00:05:12.71" />
                    <SPLIT distance="600" swimtime="00:06:17.07" />
                    <SPLIT distance="700" swimtime="00:07:21.37" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="573" eventid="15" swimtime="00:00:21.58" lane="1" heatid="15008" />
                <RESULT resultid="574" eventid="21" swimtime="00:01:51.35" reactiontime="+86" lane="1" heatid="21006">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:52.50" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="575" eventid="23" swimtime="00:03:56.92" lane="3" heatid="23001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:53.02" />
                    <SPLIT distance="200" swimtime="00:01:54.50" />
                    <SPLIT distance="300" swimtime="00:02:56.04" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY number="1" gender="M" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="532" eventid="25" swimtime="00:02:51.71" lane="5" heatid="25001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:42.66" />
                    <SPLIT distance="200" swimtime="00:01:25.21" />
                    <SPLIT distance="300" swimtime="00:02:06.46" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="195" number="1" />
                    <RELAYPOSITION athleteid="202" number="2" />
                    <RELAYPOSITION athleteid="196" number="3" />
                    <RELAYPOSITION athleteid="203" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" gender="F" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="534" eventid="24" swimtime="00:03:05.71" lane="4" heatid="24002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:48.33" />
                    <SPLIT distance="200" swimtime="00:01:33.25" />
                    <SPLIT distance="300" swimtime="00:02:17.64" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="198" number="1" />
                    <RELAYPOSITION athleteid="197" number="2" />
                    <RELAYPOSITION athleteid="201" number="3" />
                    <RELAYPOSITION athleteid="200" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" gender="X" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="720" eventid="13" swimtime="00:01:17.88" lane="4" heatid="13002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:40.10" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="197" number="1" />
                    <RELAYPOSITION athleteid="202" number="2" />
                    <RELAYPOSITION athleteid="196" number="3" />
                    <RELAYPOSITION athleteid="201" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB name="TC Marzahn e.V." nation="GER" region="21" code="0">
          <ATHLETES>
            <ATHLETE athleteid="77" birthdate="1977-01-01" gender="F" lastname="Lopez" firstname="Annett" license="0">
              <RESULTS>
                <RESULT resultid="197" eventid="1" swimtime="00:04:33.73" reactiontime="+96" lane="4" heatid="1003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:02.70" />
                    <SPLIT distance="200" swimtime="00:02:12.99" />
                    <SPLIT distance="300" swimtime="00:03:24.53" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="198" eventid="7" swimtime="00:00:56.65" reactiontime="+99" lane="6" heatid="7007" />
                <RESULT resultid="199" eventid="14" swimtime="00:00:25.34" lane="8" heatid="14008" />
                <RESULT resultid="200" eventid="20" swimtime="00:02:05.09" reactiontime="+82" lane="8" heatid="20006">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:58.81" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="78" birthdate="1971-01-01" gender="M" lastname="Tech" firstname="Matthias" license="0">
              <RESULTS>
                <RESULT resultid="201" eventid="6" swimtime="00:00:20.28" lane="5" heatid="6003" />
                <RESULT resultid="202" eventid="8" swimtime="00:00:52.16" reactiontime="+99" lane="3" heatid="8006" />
                <RESULT resultid="203" eventid="12" swimtime="00:00:25.50" lane="3" heatid="12002" />
                <RESULT resultid="204" eventid="15" swimtime="00:00:22.37" lane="5" heatid="15007" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="Tc submarin Pößneck" nation="GER" region="35" code="174116000">
          <ATHLETES>
            <ATHLETE athleteid="3" birthdate="2005-01-01" gender="F" lastname="Heinze" firstname="Charlotte" license="0">
              <RESULTS>
                <RESULT resultid="8" eventid="5" swimtime="00:00:19.04" lane="1" heatid="5004" />
                <RESULT resultid="9" eventid="7" swimtime="00:00:48.42" reactiontime="+93" lane="2" heatid="7008" />
                <RESULT resultid="10" eventid="18" swimtime="00:00:44.38" reactiontime="+97" lane="1" heatid="18004" />
                <RESULT resultid="11" eventid="22" swimtime="00:03:47.54" lane="6" heatid="22001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:52.78" />
                    <SPLIT distance="200" swimtime="00:01:49.22" />
                    <SPLIT distance="300" swimtime="00:02:49.78" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="4" birthdate="2007-01-01" gender="F" lastname="Näther" firstname="Emilia" license="0">
              <RESULTS>
                <RESULT resultid="12" eventid="1" swimtime="00:04:07.24" reactiontime="+96" lane="8" heatid="1004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:56.03" />
                    <SPLIT distance="200" swimtime="00:02:00.50" />
                    <SPLIT distance="300" swimtime="00:03:06.14" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="13" eventid="5" swimtime="00:00:19.64" lane="3" heatid="5003" />
                <RESULT resultid="14" eventid="7" swimtime="00:00:47.85" reactiontime="+95" lane="2" heatid="7009" />
                <RESULT resultid="15" eventid="14" swimtime="00:00:20.71" lane="1" heatid="14011" />
                <RESULT resultid="16" eventid="18" swimtime="00:00:48.39" reactiontime="+88" lane="6" heatid="18003" />
                <RESULT resultid="17" eventid="22" swimtime="00:04:06.51" lane="2" heatid="22001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:53.96" />
                    <SPLIT distance="200" swimtime="00:01:58.29" />
                    <SPLIT distance="300" swimtime="00:03:04.18" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="5" birthdate="2008-01-01" gender="M" lastname="Korn" firstname="Kristoph" license="0">
              <RESULTS>
                <RESULT resultid="18" eventid="6" swimtime="00:00:22.52" lane="3" heatid="6002" />
                <RESULT resultid="19" eventid="8" swimtime="00:00:57.30" reactiontime="+94" lane="8" heatid="8006" />
                <RESULT resultid="20" eventid="10" swimtime="00:08:58.63" reactiontime="+90" lane="7" heatid="10001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:00.13" />
                    <SPLIT distance="200" swimtime="00:02:17.04" />
                    <SPLIT distance="300" swimtime="00:03:35.85" />
                    <SPLIT distance="400" swimtime="00:04:59.48" />
                    <SPLIT distance="500" swimtime="00:06:17.98" />
                    <SPLIT distance="600" swimtime="00:07:14.43" />
                    <SPLIT distance="700" swimtime="00:07:43.02" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="21" eventid="15" status="DSQ" swimtime="00:00:23.96" lane="5" heatid="15005" comment="Falscher Start." />
                <RESULT resultid="22" eventid="21" swimtime="00:02:08.96" reactiontime="+77" lane="8" heatid="21005">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:59.65" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="TC Weimar" nation="GER" region="35" code="0">
          <ATHLETES>
            <ATHLETE athleteid="295" birthdate="2009-01-01" gender="M" lastname="Klabunde" firstname="Kalle" license="0">
              <RESULTS>
                <RESULT resultid="710" eventid="2" swimtime="00:04:53.04" lane="8" heatid="2003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:07.57" />
                    <SPLIT distance="200" swimtime="00:02:24.27" />
                    <SPLIT distance="300" swimtime="00:03:41.89" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="711" eventid="4" swimtime="00:00:31.44" lane="4" heatid="4001" />
                <RESULT resultid="712" eventid="8" swimtime="00:01:07.40" lane="7" heatid="8005" />
                <RESULT resultid="713" eventid="15" swimtime="00:00:27.25" lane="7" heatid="15004" />
                <RESULT resultid="714" eventid="21" swimtime="00:02:21.04" lane="6" heatid="21004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:07.30" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="296" birthdate="2011-01-01" gender="M" lastname="Bellmann" firstname="Lennart" license="0">
              <RESULTS>
                <RESULT resultid="715" eventid="2" swimtime="00:04:28.55" lane="6" heatid="2003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:04.28" />
                    <SPLIT distance="200" swimtime="00:02:14.34" />
                    <SPLIT distance="300" swimtime="00:03:23.50" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="716" eventid="8" swimtime="00:00:55.24" lane="1" heatid="8006" />
                <RESULT resultid="717" eventid="15" swimtime="00:00:24.67" lane="2" heatid="15005" />
                <RESULT resultid="718" eventid="19" swimtime="00:01:02.63" lane="6" heatid="19001" />
                <RESULT resultid="719" eventid="21" swimtime="00:02:07.38" reactiontime="+85" lane="3" heatid="21004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:02.96" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="TSC - Schwandorf e.V." nation="GER" region="34" code="0">
          <ATHLETES>
            <ATHLETE athleteid="28" birthdate="2007-01-01" gender="F" lastname="Rödl" firstname="Emily" license="0">
              <RESULTS>
                <RESULT resultid="65" eventid="1" swimtime="00:03:53.68" reactiontime="+96" lane="4" heatid="1004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:53.96" />
                    <SPLIT distance="200" swimtime="00:01:54.92" />
                    <SPLIT distance="300" swimtime="00:02:56.17" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="66" eventid="5" swimtime="00:00:20.04" lane="2" heatid="5003" />
                <RESULT resultid="67" eventid="7" swimtime="00:00:48.08" reactiontime="+75" lane="3" heatid="7008" />
                <RESULT resultid="68" eventid="18" swimtime="00:00:47.26" reactiontime="+61" lane="3" heatid="18003" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="29" birthdate="2004-01-01" gender="F" lastname="Kohler" firstname="Nina" license="0">
              <RESULTS>
                <RESULT resultid="69" eventid="5" swimtime="00:00:17.76" lane="6" heatid="5004" />
                <RESULT resultid="70" eventid="7" swimtime="00:00:44.23" reactiontime="+88" lane="2" heatid="7010" />
                <RESULT resultid="71" eventid="14" swimtime="00:00:19.87" lane="2" heatid="14011" />
                <RESULT resultid="72" eventid="18" swimtime="00:00:41.73" reactiontime="+77" lane="6" heatid="18004" />
                <RESULT resultid="73" eventid="20" swimtime="00:01:39.23" reactiontime="+90" lane="6" heatid="20007">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:48.68" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="TSC Rostock 1957 e.V." nation="GER" region="22" code="0">
          <ATHLETES>
            <ATHLETE athleteid="139" birthdate="1998-01-01" gender="F" lastname="Dethloff" firstname="Lisa" license="0">
              <RESULTS>
                <RESULT resultid="388" eventid="7" status="DNS" swimtime="00:00:00.00" lane="7" heatid="7009" />
                <RESULT resultid="389" eventid="18" swimtime="00:00:56.26" lane="4" heatid="18003" />
                <RESULT resultid="390" eventid="20" status="DNS" swimtime="00:00:00.00" lane="3" heatid="20001" />
                <RESULT resultid="391" eventid="22" status="DNS" swimtime="00:00:00.00" lane="5" heatid="22001" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
      </CLUBS>
    </MEET>
  </MEETS>
</LENEX>
