<?xml version="1.0" encoding="UTF-8"?>
<LENEX version="3.0">
  <CONSTRUCTOR name="EasyWk" version="5.23 BETA" registration="">
    <CONTACT name="Bjoern Stickan" internet="http://www.easywk.de" email="info@easywk.de" />
  </CONSTRUCTOR>
  <MEETS>
    <MEET city="Erfurt" course="LCM" name="Offene Thüringer Landesmeisterschaften im Finswimming" nation="GER" organizer="Tauchsportclub Erfurt e.V." hostclub="Tauchsportverband Thüringern e.V." deadline="2023-01-15" timing="AUTOMATIC">
      <CONTACT email="thlm@fs-ergebnisse.de" internet="www.fs-ergebnisse.de/2023/thlm" name="Delcuvé, Sabine" phone="0160 99161353" />
      <AGEDATE type="YEAR" value="2023-01-01" />
      <SESSIONS>
        <SESSION number="1" date="2023-01-21" daytime="09:20" officialmeeting="08:30" warmupfrom="08:00">
          <EVENTS>
            <EVENT eventid="1" number="1" gender="F" round="TIM">
              <SWIMSTYLE stroke="APNEA" relaycount="1" distance="50" />
              <FEE value="500" currency="EUR" />
              <HEATS>
                <HEAT heatid="1001" number="1" />
                <HEAT heatid="1002" number="2" />
                <HEAT heatid="1003" number="3" />
                <HEAT heatid="1004" number="4" />
                <HEAT heatid="1005" number="5" />
                <HEAT heatid="1006" number="6" />
                <HEAT heatid="1007" number="7" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="9" agemin="14" name="Thüringen: Kategorie G (Jg.2014 u.j.)" />
                <AGEGROUP agegroupid="2" agemax="10" agemin="14" name="Thüringen: Kategorie F (Jg.2013)" />
                <AGEGROUP agegroupid="3" agemax="11" agemin="14" name="Thüringen: Kategorie E (Jg.2012)" />
                <AGEGROUP agegroupid="4" agemax="13" agemin="14" name="Thüringen: Kategorie D (Jg.2010/2011)" />
                <AGEGROUP agegroupid="5" agemax="15" agemin="14" name="Thüringen: Kategorie C (Jg.2008/2009)">
                  <RANKINGS>
                    <RANKING place="8" resultid="505" />
                    <RANKING place="6" resultid="509" />
                    <RANKING place="4" resultid="517" />
                    <RANKING place="2" resultid="594" />
                    <RANKING place="1" resultid="765" />
                    <RANKING place="3" resultid="767" />
                    <RANKING place="7" resultid="768" />
                    <RANKING place="5" resultid="900" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6" agemax="17" agemin="16" name="Thüringen: Kategorie B (Jg.2006/2007)">
                  <RANKINGS>
                    <RANKING place="1" resultid="258" />
                    <RANKING place="4" resultid="489" />
                    <RANKING place="2" resultid="569" />
                    <RANKING place="3" resultid="766" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7" agemax="30" agemin="18" name="Thüringen: Kategorie A (Jg.2005 u.ä.)">
                  <RANKINGS>
                    <RANKING place="2" resultid="257" />
                    <RANKING place="1" resultid="338" />
                    <RANKING place="3" resultid="563" />
                    <RANKING place="4" resultid="764" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8" agemax="34" agemin="29" name="Thüringen: Master A (Jg.1989-1994)" />
                <AGEGROUP agegroupid="9" agemax="44" agemin="35" name="Thüringen: Master B (Jg.1979-1988)" />
                <AGEGROUP agegroupid="10" agemax="54" agemin="45" name="Thüringen: Master C (Jg.1969-1978)" />
                <AGEGROUP agegroupid="11" agemax="64" agemin="55" name="Thüringen: Master D (Jg.1959-1968)" />
                <AGEGROUP agegroupid="12" agemax="123" agemin="65" name="Thüringen: Master E (Jg.1958 u.ä.)" />
                <AGEGROUP agegroupid="13" agemax="123" agemin="29" name="Offene Wertung Master">
                  <RANKINGS>
                    <RANKING place="1" resultid="675" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="14" agemax="30" agemin="14" name="Offene Wertung">
                  <RANKINGS>
                    <RANKING place="2" resultid="24" />
                    <RANKING place="8" resultid="25" />
                    <RANKING place="24" resultid="26" />
                    <RANKING place="14" resultid="27" />
                    <RANKING place="41" resultid="28" />
                    <RANKING place="20" resultid="57" />
                    <RANKING place="21" resultid="91" />
                    <RANKING place="22" resultid="92" />
                    <RANKING place="28" resultid="93" />
                    <RANKING place="32" resultid="94" />
                    <RANKING place="35" resultid="95" />
                    <RANKING place="38" resultid="96" />
                    <RANKING place="36" resultid="116" />
                    <RANKING place="47" resultid="117" />
                    <RANKING place="4" resultid="128" />
                    <RANKING place="6" resultid="137" />
                    <RANKING place="12" resultid="171" />
                    <RANKING place="16" resultid="172" />
                    <RANKING place="23" resultid="173" />
                    <RANKING place="10" resultid="257" />
                    <RANKING place="13" resultid="258" />
                    <RANKING place="15" resultid="289" />
                    <RANKING place="7" resultid="338" />
                    <RANKING place="5" resultid="404" />
                    <RANKING place="19" resultid="445" />
                    <RANKING place="26" resultid="446" />
                    <RANKING place="25" resultid="447" />
                    <RANKING place="37" resultid="448" />
                    <RANKING place="33" resultid="489" />
                    <RANKING place="46" resultid="505" />
                    <RANKING place="44" resultid="509" />
                    <RANKING place="39" resultid="517" />
                    <RANKING place="40" resultid="535" />
                    <RANKING place="30" resultid="539" />
                    <RANKING place="11" resultid="563" />
                    <RANKING place="18" resultid="569" />
                    <RANKING place="27" resultid="594" />
                    <RANKING place="1" resultid="679" />
                    <RANKING place="3" resultid="683" />
                    <RANKING place="30" resultid="764" />
                    <RANKING place="17" resultid="765" />
                    <RANKING place="29" resultid="766" />
                    <RANKING place="34" resultid="767" />
                    <RANKING place="45" resultid="768" />
                    <RANKING place="9" resultid="845" />
                    <RANKING place="43" resultid="854" />
                    <RANKING place="42" resultid="900" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="2" number="2" gender="M" round="TIM">
              <SWIMSTYLE stroke="APNEA" relaycount="1" distance="50" />
              <FEE value="500" currency="EUR" />
              <HEATS>
                <HEAT heatid="2001" number="1" />
                <HEAT heatid="2002" number="2" />
                <HEAT heatid="2003" number="3" />
                <HEAT heatid="2004" number="4" />
                <HEAT heatid="2005" number="5" />
                <HEAT heatid="2006" number="6" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="9" agemin="14" name="Thüringen: Kategorie G (Jg.2014 u.j.)" />
                <AGEGROUP agegroupid="2" agemax="10" agemin="14" name="Thüringen: Kategorie F (Jg.2013)" />
                <AGEGROUP agegroupid="3" agemax="11" agemin="14" name="Thüringen: Kategorie E (Jg.2012)" />
                <AGEGROUP agegroupid="4" agemax="13" agemin="14" name="Thüringen: Kategorie D (Jg.2010/2011)" />
                <AGEGROUP agegroupid="5" agemax="15" agemin="14" name="Thüringen: Kategorie C (Jg.2008/2009)">
                  <RANKINGS>
                    <RANKING place="1" resultid="340" />
                    <RANKING place="2" resultid="501" />
                    <RANKING place="5" resultid="581" />
                    <RANKING place="3" resultid="598" />
                    <RANKING place="4" resultid="771" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6" agemax="17" agemin="16" name="Thüringen: Kategorie B (Jg.2006/2007)">
                  <RANKINGS>
                    <RANKING place="2" resultid="341" />
                    <RANKING place="1" resultid="769" />
                    <RANKING place="3" resultid="895" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7" agemax="30" agemin="18" name="Thüringen: Kategorie A (Jg.2005 u.ä.)">
                  <RANKINGS>
                    <RANKING place="2" resultid="339" />
                    <RANKING place="3" resultid="342" />
                    <RANKING place="1" resultid="878" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8" agemax="34" agemin="29" name="Thüringen: Master A (Jg.1989-1994)" />
                <AGEGROUP agegroupid="9" agemax="44" agemin="35" name="Thüringen: Master B (Jg.1979-1988)" />
                <AGEGROUP agegroupid="10" agemax="54" agemin="45" name="Thüringen: Master C (Jg.1969-1978)">
                  <RANKINGS>
                    <RANKING place="5" resultid="347" />
                    <RANKING place="2" resultid="555" />
                    <RANKING place="1" resultid="770" />
                    <RANKING place="3" resultid="772" />
                    <RANKING place="4" resultid="773" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11" agemax="64" agemin="55" name="Thüringen: Master D (Jg.1959-1968)">
                  <RANKINGS>
                    <RANKING place="1" resultid="344" />
                    <RANKING place="2" resultid="346" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="12" agemax="123" agemin="65" name="Thüringen: Master E (Jg.1958 u.ä.)">
                  <RANKINGS>
                    <RANKING place="1" resultid="345" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="13" agemax="123" agemin="28" name="Offene Wertung Master">
                  <RANKINGS>
                    <RANKING place="6" resultid="344" />
                    <RANKING place="7" resultid="345" />
                    <RANKING place="10" resultid="346" />
                    <RANKING place="9" resultid="347" />
                    <RANKING place="3" resultid="555" />
                    <RANKING place="1" resultid="770" />
                    <RANKING place="5" resultid="772" />
                    <RANKING place="8" resultid="773" />
                    <RANKING place="4" resultid="818" />
                    <RANKING place="2" resultid="821" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="14" agemax="29" agemin="14" name="Offene Wertung">
                  <RANKINGS>
                    <RANKING place="7" resultid="29" />
                    <RANKING place="17" resultid="30" />
                    <RANKING place="26" resultid="31" />
                    <RANKING place="33" resultid="41" />
                    <RANKING place="32" resultid="42" />
                    <RANKING place="1" resultid="50" />
                    <RANKING place="12" resultid="97" />
                    <RANKING place="21" resultid="98" />
                    <RANKING place="23" resultid="99" />
                    <RANKING place="31" resultid="100" />
                    <RANKING place="15" resultid="174" />
                    <RANKING place="11" resultid="175" />
                    <RANKING place="6" resultid="204" />
                    <RANKING place="16" resultid="206" />
                    <RANKING place="25" resultid="207" />
                    <RANKING place="9" resultid="339" />
                    <RANKING place="13" resultid="340" />
                    <RANKING place="20" resultid="341" />
                    <RANKING place="22" resultid="342" />
                    <RANKING place="19" resultid="405" />
                    <RANKING place="5" resultid="449" />
                    <RANKING place="14" resultid="450" />
                    <RANKING place="27" resultid="451" />
                    <RANKING place="24" resultid="501" />
                    <RANKING place="4" resultid="527" />
                    <RANKING place="10" resultid="531" />
                    <RANKING place="34" resultid="543" />
                    <RANKING place="35" resultid="581" />
                    <RANKING place="28" resultid="598" />
                    <RANKING place="2" resultid="769" />
                    <RANKING place="30" resultid="771" />
                    <RANKING place="8" resultid="832" />
                    <RANKING place="18" resultid="840" />
                    <RANKING place="3" resultid="878" />
                    <RANKING place="29" resultid="895" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="3" number="3" gender="F" round="TIM">
              <SWIMSTYLE stroke="IMMERSION" technique="DIVE" relaycount="1" distance="50" />
              <FEE value="500" currency="EUR" />
              <HEATS>
                <HEAT heatid="3001" number="1" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="9" agemin="12" name="Thüringen: Kategorie G (Jg.2014 u.j.)" />
                <AGEGROUP agegroupid="2" agemax="10" agemin="12" name="Thüringen: Kategorie F (Jg.2013)" />
                <AGEGROUP agegroupid="3" agemax="11" agemin="12" name="Thüringen: Kategorie E (Jg.2012)" />
                <AGEGROUP agegroupid="4" agemax="13" agemin="12" name="Thüringen: Kategorie D (Jg.2010/2011)">
                  <RANKINGS>
                    <RANKING place="2" resultid="277" />
                    <RANKING place="5" resultid="605" />
                    <RANKING place="1" resultid="809" />
                    <RANKING place="3" resultid="913" />
                    <RANKING place="6" resultid="919" />
                    <RANKING place="4" resultid="925" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="13" agemin="14" name="Thüringen: Kategorie C (Jg.2008/2009)" />
                <AGEGROUP agegroupid="6" agemax="13" agemin="16" name="Thüringen: Kategorie B (Jg.2006/2007)" />
                <AGEGROUP agegroupid="7" agemax="13" agemin="18" name="Thüringen: Kategorie A (Jg.2005 u.ä.)" />
                <AGEGROUP agegroupid="8" agemax="13" agemin="29" name="Thüringen: Master A (Jg.1989-1994)" />
                <AGEGROUP agegroupid="9" agemax="13" agemin="35" name="Thüringen: Master B (Jg.1979-1988)" />
                <AGEGROUP agegroupid="10" agemax="13" agemin="45" name="Thüringen: Master C (Jg.1969-1978)" />
                <AGEGROUP agegroupid="11" agemax="13" agemin="55" name="Thüringen: Master D (Jg.1959-1968)" />
                <AGEGROUP agegroupid="12" agemax="13" agemin="65" name="Thüringen: Master E (Jg.1958 u.ä.)" />
                <AGEGROUP agegroupid="13" agemax="13" agemin="29" name="Offene Wertung Master" />
                <AGEGROUP agegroupid="14" agemax="13" agemin="12" name="Offene Wertung">
                  <RANKINGS>
                    <RANKING place="2" resultid="277" />
                    <RANKING place="4" resultid="547" />
                    <RANKING place="6" resultid="605" />
                    <RANKING place="1" resultid="809" />
                    <RANKING place="3" resultid="913" />
                    <RANKING place="7" resultid="919" />
                    <RANKING place="5" resultid="925" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="4" number="4" gender="M" round="TIM">
              <SWIMSTYLE stroke="IMMERSION" technique="DIVE" relaycount="1" distance="50" />
              <FEE value="500" currency="EUR" />
              <HEATS>
                <HEAT heatid="4001" number="1" />
                <HEAT heatid="4002" number="2" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="9" agemin="12" name="Thüringen: Kategorie G (Jg.2014 u.j.)" />
                <AGEGROUP agegroupid="2" agemax="10" agemin="12" name="Thüringen: Kategorie F (Jg.2013)" />
                <AGEGROUP agegroupid="3" agemax="11" agemin="12" name="Thüringen: Kategorie E (Jg.2012)" />
                <AGEGROUP agegroupid="4" agemax="13" agemin="12" name="Thüringen: Kategorie D (Jg.2010/2011)">
                  <RANKINGS>
                    <RANKING place="7" resultid="278" />
                    <RANKING place="4" resultid="377" />
                    <RANKING place="2" resultid="378" />
                    <RANKING place="9" resultid="609" />
                    <RANKING place="6" resultid="620" />
                    <RANKING place="5" resultid="810" />
                    <RANKING place="3" resultid="811" />
                    <RANKING place="1" resultid="812" />
                    <RANKING place="8" resultid="939" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="13" agemin="14" name="Thüringen: Kategorie C (Jg.2008/2009)" />
                <AGEGROUP agegroupid="6" agemax="13" agemin="16" name="Thüringen: Kategorie B (Jg.2006/2007)" />
                <AGEGROUP agegroupid="7" agemax="13" agemin="18" name="Thüringen: Kategorie A (Jg.2005 u.ä.)" />
                <AGEGROUP agegroupid="8" agemax="13" agemin="29" name="Thüringen: Master A (Jg.1989-1994)" />
                <AGEGROUP agegroupid="9" agemax="13" agemin="35" name="Thüringen: Master B (Jg.1979-1988)" />
                <AGEGROUP agegroupid="10" agemax="13" agemin="45" name="Thüringen: Master C (Jg.1969-1978)" />
                <AGEGROUP agegroupid="11" agemax="13" agemin="55" name="Thüringen: Master D (Jg.1959-1968)" />
                <AGEGROUP agegroupid="12" agemax="13" agemin="65" name="Thüringen: Master E (Jg.1958 u.ä.)" />
                <AGEGROUP agegroupid="13" agemax="13" agemin="28" name="Offene Wertung Master" />
                <AGEGROUP agegroupid="14" agemax="13" agemin="12" name="Offene Wertung">
                  <RANKINGS>
                    <RANKING place="2" resultid="111" />
                    <RANKING place="8" resultid="278" />
                    <RANKING place="5" resultid="377" />
                    <RANKING place="3" resultid="378" />
                    <RANKING place="10" resultid="609" />
                    <RANKING place="7" resultid="620" />
                    <RANKING place="6" resultid="810" />
                    <RANKING place="4" resultid="811" />
                    <RANKING place="1" resultid="812" />
                    <RANKING place="9" resultid="939" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="5" number="5" gender="F" round="TIM">
              <SWIMSTYLE stroke="FLY" technique="KICK" relaycount="1" distance="50" />
              <FEE value="500" currency="EUR" />
              <HEATS>
                <HEAT heatid="5001" number="1" />
                <HEAT heatid="5002" number="2" />
                <HEAT heatid="5003" number="3" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="9" agemin="1" name="Thüringen: Kategorie G (Jg.2014 u.j.)">
                  <RANKINGS>
                    <RANKING place="2" resultid="523" />
                    <RANKING place="1" resultid="952" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2" agemax="10" agemin="10" name="Thüringen: Kategorie F (Jg.2013)">
                  <RANKINGS>
                    <RANKING place="4" resultid="259" />
                    <RANKING place="1" resultid="261" />
                    <RANKING place="2" resultid="640" />
                    <RANKING place="3" resultid="774" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3" agemax="11" agemin="11" name="Thüringen: Kategorie E (Jg.2012)">
                  <RANKINGS>
                    <RANKING place="1" resultid="260" />
                    <RANKING place="7" resultid="348" />
                    <RANKING place="5" resultid="349" />
                    <RANKING place="4" resultid="351" />
                    <RANKING place="6" resultid="775" />
                    <RANKING place="3" resultid="776" />
                    <RANKING place="2" resultid="947" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="11" agemin="12" name="Thüringen: Kategorie D (Jg.2010/2011)" />
                <AGEGROUP agegroupid="5" agemax="11" agemin="14" name="Thüringen: Kategorie C (Jg.2008/2009)" />
                <AGEGROUP agegroupid="6" agemax="11" agemin="16" name="Thüringen: Kategorie B (Jg.2006/2007)" />
                <AGEGROUP agegroupid="7" agemax="11" agemin="18" name="Thüringen: Kategorie A (Jg.2005 u.ä.)" />
                <AGEGROUP agegroupid="8" agemax="11" agemin="29" name="Thüringen: Master A (Jg.1989-1994)" />
                <AGEGROUP agegroupid="9" agemax="11" agemin="35" name="Thüringen: Master B (Jg.1979-1988)" />
                <AGEGROUP agegroupid="10" agemax="11" agemin="45" name="Thüringen: Master C (Jg.1969-1978)" />
                <AGEGROUP agegroupid="11" agemax="11" agemin="55" name="Thüringen: Master D (Jg.1959-1968)" />
                <AGEGROUP agegroupid="12" agemax="11" agemin="65" name="Thüringen: Master E (Jg.1958 u.ä.)" />
                <AGEGROUP agegroupid="13" agemax="11" agemin="29" name="Offene Wertung Master" />
                <AGEGROUP agegroupid="14" agemax="11" agemin="1" name="Offene Wertung">
                  <RANKINGS>
                    <RANKING place="5" resultid="176" />
                    <RANKING place="8" resultid="177" />
                    <RANKING place="16" resultid="259" />
                    <RANKING place="1" resultid="260" />
                    <RANKING place="10" resultid="261" />
                    <RANKING place="12" resultid="290" />
                    <RANKING place="13" resultid="348" />
                    <RANKING place="9" resultid="349" />
                    <RANKING place="7" resultid="351" />
                    <RANKING place="6" resultid="452" />
                    <RANKING place="4" resultid="453" />
                    <RANKING place="18" resultid="523" />
                    <RANKING place="14" resultid="640" />
                    <RANKING place="15" resultid="774" />
                    <RANKING place="11" resultid="775" />
                    <RANKING place="3" resultid="776" />
                    <RANKING place="2" resultid="947" />
                    <RANKING place="17" resultid="952" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="6" number="6" gender="M" round="TIM">
              <SWIMSTYLE stroke="FLY" technique="KICK" relaycount="1" distance="50" />
              <FEE value="500" currency="EUR" />
              <HEATS>
                <HEAT heatid="6001" number="1" />
                <HEAT heatid="6002" number="2" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="9" agemin="1" name="Thüringen: Kategorie G (Jg.2014 u.j.)">
                  <RANKINGS>
                    <RANKING place="1" resultid="655" />
                    <RANKING place="2" resultid="664" />
                    <RANKING place="3" resultid="672" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2" agemax="10" agemin="10" name="Thüringen: Kategorie F (Jg.2013)" />
                <AGEGROUP agegroupid="3" agemax="11" agemin="11" name="Thüringen: Kategorie E (Jg.2012)">
                  <RANKINGS>
                    <RANKING place="1" resultid="635" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="11" agemin="12" name="Thüringen: Kategorie D (Jg.2010/2011)" />
                <AGEGROUP agegroupid="5" agemax="11" agemin="14" name="Thüringen: Kategorie C (Jg.2008/2009)" />
                <AGEGROUP agegroupid="6" agemax="11" agemin="16" name="Thüringen: Kategorie B (Jg.2006/2007)" />
                <AGEGROUP agegroupid="7" agemax="11" agemin="18" name="Thüringen: Kategorie A (Jg.2005 u.ä.)" />
                <AGEGROUP agegroupid="8" agemax="11" agemin="29" name="Thüringen: Master A (Jg.1989-1994)" />
                <AGEGROUP agegroupid="9" agemax="11" agemin="35" name="Thüringen: Master B (Jg.1979-1988)" />
                <AGEGROUP agegroupid="10" agemax="11" agemin="45" name="Thüringen: Master C (Jg.1969-1978)" />
                <AGEGROUP agegroupid="11" agemax="11" agemin="55" name="Thüringen: Master D (Jg.1959-1968)" />
                <AGEGROUP agegroupid="12" agemax="11" agemin="65" name="Thüringen: Master E (Jg.1958 u.ä.)" />
                <AGEGROUP agegroupid="13" agemax="11" agemin="28" name="Offene Wertung Master" />
                <AGEGROUP agegroupid="14" agemax="11" agemin="1" name="Offene Wertung">
                  <RANKINGS>
                    <RANKING place="2" resultid="454" />
                    <RANKING place="3" resultid="455" />
                    <RANKING place="1" resultid="635" />
                    <RANKING place="4" resultid="655" />
                    <RANKING place="5" resultid="664" />
                    <RANKING place="6" resultid="672" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="7" number="7" gender="X" round="TIM">
              <SWIMSTYLE stroke="SURFACE" relaycount="1" distance="800" />
              <FEE value="500" currency="EUR" />
              <HEATS>
                <HEAT heatid="7001" number="1" />
                <HEAT heatid="7002" number="2" />
                <HEAT heatid="7003" number="3" />
                <HEAT heatid="7004" number="4" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="9" agemin="11" name="weiblich Thüringen: Kategorie G (Jg.2014 u.j.)" />
                <AGEGROUP agegroupid="2" agemax="10" agemin="11" name="weiblich Thüringen: Kategorie F (Jg.2013)" />
                <AGEGROUP agegroupid="3" agemax="11" agemin="11" name="weiblich Thüringen: Kategorie E (Jg.2012)" />
                <AGEGROUP agegroupid="4" agemax="13" agemin="12" name="weiblich Thüringen: Kategorie D (Jg.2010/2011)" />
                <AGEGROUP agegroupid="5" agemax="15" agemin="14" name="weiblich Thüringen: Kategorie C (Jg.2008/2009)">
                  <RANKINGS>
                    <RANKING place="1" resultid="813" />
                    <RANKING place="2" resultid="901" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6" agemax="17" agemin="16" name="weiblich Thüringen: Kategorie B (Jg.2006/2007)">
                  <RANKINGS>
                    <RANKING place="1" resultid="490" />
                    <RANKING place="2" resultid="494" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7" agemax="30" agemin="18" name="weiblich Thüringen: Kategorie A (Jg.2005 u.ä.)">
                  <RANKINGS>
                    <RANKING place="2" resultid="474" />
                    <RANKING place="1" resultid="478" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8" agemax="34" agemin="29" name="weiblich Thüringen: Master A (Jg.1989-1994)" />
                <AGEGROUP agegroupid="9" agemax="44" agemin="35" name="weiblich Thüringen: Master B (Jg.1979-1988)" />
                <AGEGROUP agegroupid="10" agemax="54" agemin="45" name="weiblich Thüringen: Master C (Jg.1969-1978)" />
                <AGEGROUP agegroupid="11" agemax="64" agemin="55" name="weiblich Thüringen: Master D (Jg.1959-1968)" />
                <AGEGROUP agegroupid="12" agemax="123" agemin="65" name="weiblich Thüringen: Master E (Jg.1958 u.ä.)" />
                <AGEGROUP agegroupid="13" agemax="123" agemin="29" name="weiblich: Offene Wertung Master" />
                <AGEGROUP agegroupid="14" agemax="30" agemin="11" name="weiblich: Offene Wertung">
                  <RANKINGS>
                    <RANKING place="5" resultid="58" />
                    <RANKING place="6" resultid="133" />
                    <RANKING place="4" resultid="188" />
                    <RANKING place="2" resultid="189" />
                    <RANKING place="10" resultid="191" />
                    <RANKING place="8" resultid="215" />
                    <RANKING place="1" resultid="413" />
                    <RANKING place="12" resultid="470" />
                    <RANKING place="11" resultid="474" />
                    <RANKING place="7" resultid="478" />
                    <RANKING place="13" resultid="490" />
                    <RANKING place="16" resultid="494" />
                    <RANKING place="9" resultid="813" />
                    <RANKING place="15" resultid="859" />
                    <RANKING place="14" resultid="901" />
                    <RANKING place="3" resultid="955" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15" agemax="9" agemin="11" name="männlich Thüringen: Kategorie G (Jg.2014 u.j.)" />
                <AGEGROUP agegroupid="16" agemax="10" agemin="11" name="männlich Thüringen: Kategorie F (Jg.2013)" />
                <AGEGROUP agegroupid="17" agemax="11" agemin="11" name="männlich Thüringen: Kategorie E (Jg.2012)" />
                <AGEGROUP agegroupid="18" agemax="13" agemin="12" name="männlich Thüringen: Kategorie D (Jg.2010/2011)" />
                <AGEGROUP agegroupid="19" agemax="15" agemin="14" name="männlich Thüringen: Kategorie C (Jg.2008/2009)">
                  <RANKINGS>
                    <RANKING place="1" resultid="814" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="20" agemax="17" agemin="16" name="männlich Thüringen: Kategorie B (Jg.2006/2007)">
                  <RANKINGS>
                    <RANKING place="1" resultid="896" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="21" agemax="30" agemin="18" name="männlich Thüringen: Kategorie A (Jg.2005 u.ä.)">
                  <RANKINGS>
                    <RANKING place="2" resultid="875" />
                    <RANKING place="1" resultid="883" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="22" agemax="34" agemin="29" name="männlich Thüringen: Master A (Jg.1989-1994)" />
                <AGEGROUP agegroupid="23" agemax="44" agemin="35" name="männlich Thüringen: Master B (Jg.1979-1988)" />
                <AGEGROUP agegroupid="24" agemax="54" agemin="45" name="männlich Thüringen: Master C (Jg.1969-1978)" />
                <AGEGROUP agegroupid="25" agemax="64" agemin="55" name="männlich Thüringen: Master D (Jg.1959-1968)" />
                <AGEGROUP agegroupid="26" agemax="123" agemin="65" name="männlich Thüringen: Master E (Jg.1958 u.ä.)" />
                <AGEGROUP agegroupid="27" agemax="123" agemin="28" name="männlich: Offene Wertung Master" />
                <AGEGROUP agegroupid="28" agemax="29" agemin="11" name="männlich: Offene Wertung">
                  <RANKINGS>
                    <RANKING place="6" resultid="46" />
                    <RANKING place="4" resultid="112" />
                    <RANKING place="1" resultid="528" />
                    <RANKING place="7" resultid="814" />
                    <RANKING place="3" resultid="875" />
                    <RANKING place="2" resultid="883" />
                    <RANKING place="5" resultid="896" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="8" number="8" gender="F" round="TIM">
              <SWIMSTYLE stroke="SURFACE" relaycount="1" distance="100" />
              <FEE value="500" currency="EUR" />
              <HEATS>
                <HEAT heatid="8001" number="1" />
                <HEAT heatid="8002" number="2" />
                <HEAT heatid="8003" number="3" />
                <HEAT heatid="8004" number="4" />
                <HEAT heatid="8005" number="5" />
                <HEAT heatid="8006" number="6" />
                <HEAT heatid="8007" number="7" />
                <HEAT heatid="8008" number="8" />
                <HEAT heatid="8009" number="9" />
                <HEAT heatid="8010" number="10" />
                <HEAT heatid="8011" number="11" />
                <HEAT heatid="8012" number="12" />
                <HEAT heatid="8013" number="13" />
                <HEAT heatid="8014" number="14" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="9" agemin="1" name="Thüringen: Kategorie G (Jg.2014 u.j.)">
                  <RANKINGS>
                    <RANKING place="3" resultid="524" />
                    <RANKING place="6" resultid="650" />
                    <RANKING place="5" resultid="652" />
                    <RANKING place="4" resultid="662" />
                    <RANKING place="1" resultid="669" />
                    <RANKING place="2" resultid="953" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2" agemax="10" agemin="10" name="Thüringen: Kategorie F (Jg.2013)">
                  <RANKINGS>
                    <RANKING place="1" resultid="221" />
                    <RANKING place="6" resultid="223" />
                    <RANKING place="3" resultid="224" />
                    <RANKING place="2" resultid="225" />
                    <RANKING place="4" resultid="296" />
                    <RANKING place="5" resultid="641" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3" agemax="11" agemin="11" name="Thüringen: Kategorie E (Jg.2012)">
                  <RANKINGS>
                    <RANKING place="1" resultid="218" />
                    <RANKING place="5" resultid="294" />
                    <RANKING place="7" resultid="295" />
                    <RANKING place="2" resultid="704" />
                    <RANKING place="3" resultid="705" />
                    <RANKING place="6" resultid="707" />
                    <RANKING place="4" resultid="948" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="13" agemin="12" name="Thüringen: Kategorie D (Jg.2010/2011)">
                  <RANKINGS>
                    <RANKING place="2" resultid="217" />
                    <RANKING place="7" resultid="219" />
                    <RANKING place="14" resultid="220" />
                    <RANKING place="3" resultid="298" />
                    <RANKING place="9" resultid="299" />
                    <RANKING place="4" resultid="300" />
                    <RANKING place="12" resultid="606" />
                    <RANKING place="10" resultid="624" />
                    <RANKING place="13" resultid="691" />
                    <RANKING place="1" resultid="693" />
                    <RANKING place="5" resultid="702" />
                    <RANKING place="16" resultid="706" />
                    <RANKING place="6" resultid="914" />
                    <RANKING place="11" resultid="920" />
                    <RANKING place="8" resultid="926" />
                    <RANKING place="15" resultid="935" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="15" agemin="14" name="Thüringen: Kategorie C (Jg.2008/2009)">
                  <RANKINGS>
                    <RANKING place="6" resultid="506" />
                    <RANKING place="4" resultid="510" />
                    <RANKING place="7" resultid="513" />
                    <RANKING place="1" resultid="595" />
                    <RANKING place="2" resultid="694" />
                    <RANKING place="3" resultid="701" />
                    <RANKING place="5" resultid="907" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6" agemax="17" agemin="16" name="Thüringen: Kategorie B (Jg.2006/2007)">
                  <RANKINGS>
                    <RANKING place="2" resultid="216" />
                    <RANKING place="1" resultid="570" />
                    <RANKING place="3" resultid="698" />
                    <RANKING place="4" resultid="699" />
                    <RANKING place="5" resultid="890" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7" agemax="30" agemin="18" name="Thüringen: Kategorie A (Jg.2005 u.ä.)">
                  <RANKINGS>
                    <RANKING place="1" resultid="564" />
                    <RANKING place="2" resultid="692" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8" agemax="34" agemin="29" name="Thüringen: Master A (Jg.1989-1994)" />
                <AGEGROUP agegroupid="9" agemax="44" agemin="35" name="Thüringen: Master B (Jg.1979-1988)">
                  <RANKINGS>
                    <RANKING place="1" resultid="696" />
                    <RANKING place="2" resultid="697" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10" agemax="54" agemin="45" name="Thüringen: Master C (Jg.1969-1978)" />
                <AGEGROUP agegroupid="11" agemax="64" agemin="55" name="Thüringen: Master D (Jg.1959-1968)">
                  <RANKINGS>
                    <RANKING place="1" resultid="703" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="12" agemax="123" agemin="65" name="Thüringen: Master E (Jg.1958 u.ä.)" />
                <AGEGROUP agegroupid="13" agemax="123" agemin="29" name="Offene Wertung Master">
                  <RANKINGS>
                    <RANKING place="3" resultid="676" />
                    <RANKING place="2" resultid="696" />
                    <RANKING place="4" resultid="697" />
                    <RANKING place="6" resultid="703" />
                    <RANKING place="1" resultid="824" />
                    <RANKING place="5" resultid="827" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="14" agemax="30" agemin="1" name="Offene Wertung">
                  <RANKINGS>
                    <RANKING place="8" resultid="1" />
                    <RANKING place="3" resultid="2" />
                    <RANKING place="11" resultid="3" />
                    <RANKING place="36" resultid="4" />
                    <RANKING place="42" resultid="5" />
                    <RANKING place="44" resultid="6" />
                    <RANKING place="15" resultid="52" />
                    <RANKING place="14" resultid="59" />
                    <RANKING place="20" resultid="60" />
                    <RANKING place="34" resultid="61" />
                    <RANKING place="26" resultid="62" />
                    <RANKING place="41" resultid="63" />
                    <RANKING place="37" resultid="64" />
                    <RANKING place="56" resultid="113" />
                    <RANKING place="44" resultid="121" />
                    <RANKING place="61" resultid="123" />
                    <RANKING place="24" resultid="134" />
                    <RANKING place="4" resultid="140" />
                    <RANKING place="6" resultid="141" />
                    <RANKING place="18" resultid="142" />
                    <RANKING place="79" resultid="143" />
                    <RANKING place="89" resultid="144" />
                    <RANKING place="94" resultid="145" />
                    <RANKING place="35" resultid="192" />
                    <RANKING place="19" resultid="216" />
                    <RANKING place="47" resultid="217" />
                    <RANKING place="50" resultid="218" />
                    <RANKING place="58" resultid="219" />
                    <RANKING place="76" resultid="220" />
                    <RANKING place="65" resultid="221" />
                    <RANKING place="88" resultid="223" />
                    <RANKING place="75" resultid="224" />
                    <RANKING place="71" resultid="225" />
                    <RANKING place="10" resultid="279" />
                    <RANKING place="9" resultid="280" />
                    <RANKING place="72" resultid="281" />
                    <RANKING place="82" resultid="282" />
                    <RANKING place="83" resultid="294" />
                    <RANKING place="93" resultid="295" />
                    <RANKING place="85" resultid="296" />
                    <RANKING place="51" resultid="298" />
                    <RANKING place="60" resultid="299" />
                    <RANKING place="52" resultid="300" />
                    <RANKING place="5" resultid="379" />
                    <RANKING place="17" resultid="380" />
                    <RANKING place="12" resultid="414" />
                    <RANKING place="23" resultid="415" />
                    <RANKING place="68" resultid="416" />
                    <RANKING place="84" resultid="417" />
                    <RANKING place="78" resultid="418" />
                    <RANKING place="80" resultid="419" />
                    <RANKING place="53" resultid="506" />
                    <RANKING place="43" resultid="510" />
                    <RANKING place="64" resultid="513" />
                    <RANKING place="92" resultid="524" />
                    <RANKING place="33" resultid="536" />
                    <RANKING place="25" resultid="540" />
                    <RANKING place="38" resultid="548" />
                    <RANKING place="48" resultid="552" />
                    <RANKING place="7" resultid="564" />
                    <RANKING place="16" resultid="570" />
                    <RANKING place="31" resultid="595" />
                    <RANKING place="73" resultid="606" />
                    <RANKING place="62" resultid="624" />
                    <RANKING place="87" resultid="641" />
                    <RANKING place="97" resultid="650" />
                    <RANKING place="96" resultid="652" />
                    <RANKING place="95" resultid="662" />
                    <RANKING place="90" resultid="669" />
                    <RANKING place="1" resultid="680" />
                    <RANKING place="2" resultid="684" />
                    <RANKING place="74" resultid="691" />
                    <RANKING place="21" resultid="692" />
                    <RANKING place="28" resultid="693" />
                    <RANKING place="32" resultid="694" />
                    <RANKING place="30" resultid="698" />
                    <RANKING place="57" resultid="699" />
                    <RANKING place="39" resultid="701" />
                    <RANKING place="54" resultid="702" />
                    <RANKING place="63" resultid="704" />
                    <RANKING place="66" resultid="705" />
                    <RANKING place="81" resultid="706" />
                    <RANKING place="86" resultid="707" />
                    <RANKING place="13" resultid="846" />
                    <RANKING place="22" resultid="849" />
                    <RANKING place="46" resultid="855" />
                    <RANKING place="27" resultid="860" />
                    <RANKING place="29" resultid="864" />
                    <RANKING place="40" resultid="868" />
                    <RANKING place="67" resultid="890" />
                    <RANKING place="49" resultid="907" />
                    <RANKING place="55" resultid="914" />
                    <RANKING place="70" resultid="920" />
                    <RANKING place="59" resultid="926" />
                    <RANKING place="77" resultid="935" />
                    <RANKING place="69" resultid="948" />
                    <RANKING place="91" resultid="953" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="9" number="9" gender="M" round="TIM">
              <SWIMSTYLE stroke="SURFACE" relaycount="1" distance="100" />
              <FEE value="500" currency="EUR" />
              <HEATS>
                <HEAT heatid="9001" number="1" />
                <HEAT heatid="9002" number="2" />
                <HEAT heatid="9003" number="3" />
                <HEAT heatid="9004" number="4" />
                <HEAT heatid="9005" number="5" />
                <HEAT heatid="9006" number="6" />
                <HEAT heatid="9007" number="7" />
                <HEAT heatid="9008" number="8" />
                <HEAT heatid="9009" number="9" />
                <HEAT heatid="9010" number="10" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="9" agemin="1" name="Thüringen: Kategorie G (Jg.2014 u.j.)">
                  <RANKINGS>
                    <RANKING place="2" resultid="302" />
                    <RANKING place="1" resultid="656" />
                    <RANKING place="4" resultid="660" />
                    <RANKING place="3" resultid="673" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2" agemax="10" agemin="10" name="Thüringen: Kategorie F (Jg.2013)">
                  <RANKINGS>
                    <RANKING place="3" resultid="226" />
                    <RANKING place="1" resultid="229" />
                    <RANKING place="2" resultid="644" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3" agemax="11" agemin="11" name="Thüringen: Kategorie E (Jg.2012)">
                  <RANKINGS>
                    <RANKING place="1" resultid="636" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="13" agemin="12" name="Thüringen: Kategorie D (Jg.2010/2011)">
                  <RANKINGS>
                    <RANKING place="8" resultid="227" />
                    <RANKING place="7" resultid="228" />
                    <RANKING place="2" resultid="310" />
                    <RANKING place="3" resultid="311" />
                    <RANKING place="9" resultid="610" />
                    <RANKING place="6" resultid="621" />
                    <RANKING place="1" resultid="711" />
                    <RANKING place="4" resultid="713" />
                    <RANKING place="5" resultid="715" />
                    <RANKING place="10" resultid="717" />
                    <RANKING place="12" resultid="931" />
                    <RANKING place="11" resultid="940" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="15" agemin="14" name="Thüringen: Kategorie C (Jg.2008/2009)">
                  <RANKINGS>
                    <RANKING place="2" resultid="308" />
                    <RANKING place="7" resultid="312" />
                    <RANKING place="5" resultid="577" />
                    <RANKING place="6" resultid="582" />
                    <RANKING place="1" resultid="586" />
                    <RANKING place="4" resultid="599" />
                    <RANKING place="3" resultid="710" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6" agemax="17" agemin="16" name="Thüringen: Kategorie B (Jg.2006/2007)">
                  <RANKINGS>
                    <RANKING place="2" resultid="306" />
                    <RANKING place="1" resultid="708" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7" agemax="30" agemin="18" name="Thüringen: Kategorie A (Jg.2005 u.ä.)">
                  <RANKINGS>
                    <RANKING place="2" resultid="305" />
                    <RANKING place="4" resultid="307" />
                    <RANKING place="1" resultid="879" />
                    <RANKING place="3" resultid="884" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8" agemax="34" agemin="29" name="Thüringen: Master A (Jg.1989-1994)" />
                <AGEGROUP agegroupid="9" agemax="44" agemin="35" name="Thüringen: Master B (Jg.1979-1988)" />
                <AGEGROUP agegroupid="10" agemax="54" agemin="45" name="Thüringen: Master C (Jg.1969-1978)">
                  <RANKINGS>
                    <RANKING place="2" resultid="556" />
                    <RANKING place="1" resultid="709" />
                    <RANKING place="3" resultid="712" />
                    <RANKING place="4" resultid="714" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11" agemax="64" agemin="55" name="Thüringen: Master D (Jg.1959-1968)" />
                <AGEGROUP agegroupid="12" agemax="123" agemin="65" name="Thüringen: Master E (Jg.1958 u.ä.)">
                  <RANKINGS>
                    <RANKING place="1" resultid="313" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="13" agemax="123" agemin="28" name="Offene Wertung Master">
                  <RANKINGS>
                    <RANKING place="6" resultid="313" />
                    <RANKING place="3" resultid="556" />
                    <RANKING place="2" resultid="709" />
                    <RANKING place="4" resultid="712" />
                    <RANKING place="7" resultid="714" />
                    <RANKING place="5" resultid="819" />
                    <RANKING place="1" resultid="957" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="14" agemax="29" agemin="1" name="Offene Wertung">
                  <RANKINGS>
                    <RANKING place="16" resultid="7" />
                    <RANKING place="24" resultid="8" />
                    <RANKING place="29" resultid="36" />
                    <RANKING place="31" resultid="37" />
                    <RANKING place="4" resultid="48" />
                    <RANKING place="15" resultid="65" />
                    <RANKING place="25" resultid="67" />
                    <RANKING place="32" resultid="68" />
                    <RANKING place="9" resultid="146" />
                    <RANKING place="7" resultid="147" />
                    <RANKING place="13" resultid="148" />
                    <RANKING place="21" resultid="193" />
                    <RANKING place="23" resultid="194" />
                    <RANKING place="54" resultid="226" />
                    <RANKING place="46" resultid="227" />
                    <RANKING place="43" resultid="228" />
                    <RANKING place="50" resultid="229" />
                    <RANKING place="55" resultid="302" />
                    <RANKING place="8" resultid="305" />
                    <RANKING place="17" resultid="306" />
                    <RANKING place="18" resultid="307" />
                    <RANKING place="19" resultid="308" />
                    <RANKING place="33" resultid="310" />
                    <RANKING place="35" resultid="311" />
                    <RANKING place="39" resultid="312" />
                    <RANKING place="1" resultid="382" />
                    <RANKING place="2" resultid="383" />
                    <RANKING place="5" resultid="384" />
                    <RANKING place="20" resultid="385" />
                    <RANKING place="22" resultid="386" />
                    <RANKING place="42" resultid="421" />
                    <RANKING place="41" resultid="422" />
                    <RANKING place="44" resultid="424" />
                    <RANKING place="28" resultid="544" />
                    <RANKING place="34" resultid="577" />
                    <RANKING place="37" resultid="582" />
                    <RANKING place="11" resultid="586" />
                    <RANKING place="27" resultid="599" />
                    <RANKING place="47" resultid="610" />
                    <RANKING place="40" resultid="621" />
                    <RANKING place="45" resultid="636" />
                    <RANKING place="51" resultid="644" />
                    <RANKING place="52" resultid="656" />
                    <RANKING place="57" resultid="660" />
                    <RANKING place="56" resultid="673" />
                    <RANKING place="3" resultid="708" />
                    <RANKING place="26" resultid="710" />
                    <RANKING place="30" resultid="711" />
                    <RANKING place="36" resultid="713" />
                    <RANKING place="38" resultid="715" />
                    <RANKING place="48" resultid="717" />
                    <RANKING place="10" resultid="833" />
                    <RANKING place="14" resultid="841" />
                    <RANKING place="6" resultid="879" />
                    <RANKING place="12" resultid="884" />
                    <RANKING place="53" resultid="931" />
                    <RANKING place="49" resultid="940" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="10" number="10" gender="X" round="TIM">
              <SWIMSTYLE stroke="IMMERSION" technique="DIVE" relaycount="1" distance="400" />
              <FEE value="500" currency="EUR" />
              <HEATS>
                <HEAT heatid="10001" number="1" />
                <HEAT heatid="10002" number="2" />
                <HEAT heatid="10003" number="3" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="9" agemin="12" name="weiblich Thüringen: Kategorie G (Jg.2014 u.j.)" />
                <AGEGROUP agegroupid="2" agemax="10" agemin="12" name="weiblich Thüringen: Kategorie F (Jg.2013)" />
                <AGEGROUP agegroupid="3" agemax="11" agemin="12" name="weiblich Thüringen: Kategorie E (Jg.2012)" />
                <AGEGROUP agegroupid="4" agemax="13" agemin="12" name="weiblich Thüringen: Kategorie D (Jg.2010/2011)" />
                <AGEGROUP agegroupid="5" agemax="15" agemin="14" name="weiblich Thüringen: Kategorie C (Jg.2008/2009)">
                  <RANKINGS>
                    <RANKING place="1" resultid="590" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6" agemax="17" agemin="16" name="weiblich Thüringen: Kategorie B (Jg.2006/2007)">
                  <RANKINGS>
                    <RANKING place="2" resultid="495" />
                    <RANKING place="1" resultid="571" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7" agemax="30" agemin="18" name="weiblich Thüringen: Kategorie A (Jg.2005 u.ä.)">
                  <RANKINGS>
                    <RANKING place="1" resultid="251" />
                    <RANKING place="3" resultid="332" />
                    <RANKING place="4" resultid="475" />
                    <RANKING place="2" resultid="479" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8" agemax="34" agemin="29" name="weiblich Thüringen: Master A (Jg.1989-1994)" />
                <AGEGROUP agegroupid="9" agemax="44" agemin="35" name="weiblich Thüringen: Master B (Jg.1979-1988)" />
                <AGEGROUP agegroupid="10" agemax="54" agemin="45" name="weiblich Thüringen: Master C (Jg.1969-1978)" />
                <AGEGROUP agegroupid="11" agemax="64" agemin="55" name="weiblich Thüringen: Master D (Jg.1959-1968)" />
                <AGEGROUP agegroupid="12" agemax="123" agemin="65" name="weiblich Thüringen: Master E (Jg.1958 u.ä.)" />
                <AGEGROUP agegroupid="13" agemax="123" agemin="29" name="weiblich: Offene Wertung Master" />
                <AGEGROUP agegroupid="14" agemax="30" agemin="12" name="weiblich: Offene Wertung">
                  <RANKINGS>
                    <RANKING place="3" resultid="55" />
                    <RANKING place="2" resultid="56" />
                    <RANKING place="1" resultid="168" />
                    <RANKING place="7" resultid="202" />
                    <RANKING place="4" resultid="251" />
                    <RANKING place="6" resultid="332" />
                    <RANKING place="9" resultid="475" />
                    <RANKING place="5" resultid="479" />
                    <RANKING place="11" resultid="495" />
                    <RANKING place="8" resultid="571" />
                    <RANKING place="10" resultid="590" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15" agemax="9" agemin="12" name="männlich Thüringen: Kategorie G (Jg.2014 u.j.)" />
                <AGEGROUP agegroupid="16" agemax="10" agemin="12" name="männlich Thüringen: Kategorie F (Jg.2013)" />
                <AGEGROUP agegroupid="17" agemax="11" agemin="12" name="männlich Thüringen: Kategorie E (Jg.2012)" />
                <AGEGROUP agegroupid="18" agemax="13" agemin="12" name="männlich Thüringen: Kategorie D (Jg.2010/2011)" />
                <AGEGROUP agegroupid="19" agemax="15" agemin="14" name="männlich Thüringen: Kategorie C (Jg.2008/2009)" />
                <AGEGROUP agegroupid="20" agemax="17" agemin="16" name="männlich Thüringen: Kategorie B (Jg.2006/2007)">
                  <RANKINGS>
                    <RANKING place="1" resultid="897" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="21" agemax="44" agemin="18" name="männlich Thüringen: Kategorie A (Jg.2005 u.ä.)">
                  <RANKINGS>
                    <RANKING place="1" resultid="331" />
                    <RANKING place="3" resultid="471" />
                    <RANKING place="2" resultid="876" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="22" agemax="34" agemin="29" name="männlich Thüringen: Master A (Jg.1989-1994)" />
                <AGEGROUP agegroupid="23" agemax="43" agemin="35" name="männlich Thüringen: Master B (Jg.1979-1988)" />
                <AGEGROUP agegroupid="24" agemax="54" agemin="45" name="männlich Thüringen: Master C (Jg.1969-1978)" />
                <AGEGROUP agegroupid="25" agemax="64" agemin="55" name="männlich Thüringen: Master D (Jg.1959-1968)" />
                <AGEGROUP agegroupid="26" agemax="123" agemin="65" name="männlich Thüringen: Master E (Jg.1958 u.ä.)" />
                <AGEGROUP agegroupid="27" agemax="123" agemin="45" name="männlich: Offene Wertung Master" />
                <AGEGROUP agegroupid="28" agemax="44" agemin="12" name="männlich: Offene Wertung">
                  <RANKINGS>
                    <RANKING place="2" resultid="22" />
                    <RANKING place="1" resultid="201" />
                    <RANKING place="3" resultid="331" />
                    <RANKING place="6" resultid="471" />
                    <RANKING place="4" resultid="876" />
                    <RANKING place="5" resultid="897" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="11" number="11" gender="F" round="TIM">
              <SWIMSTYLE stroke="SURFACE" relaycount="1" distance="50" />
              <FEE value="500" currency="EUR" />
              <HEATS>
                <HEAT heatid="11001" number="1" />
                <HEAT heatid="11002" number="2" />
                <HEAT heatid="11003" number="3" />
                <HEAT heatid="11004" number="4" />
                <HEAT heatid="11005" number="5" />
                <HEAT heatid="11006" number="6" />
                <HEAT heatid="11007" number="7" />
                <HEAT heatid="11008" number="8" />
                <HEAT heatid="11009" number="9" />
                <HEAT heatid="11010" number="10" />
                <HEAT heatid="11011" number="11" />
                <HEAT heatid="11012" number="12" />
                <HEAT heatid="11013" number="13" />
                <HEAT heatid="11014" number="14" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="9" agemin="1" name="Thüringen: Kategorie G (Jg.2014 u.j.)">
                  <RANKINGS>
                    <RANKING place="6" resultid="272" />
                    <RANKING place="7" resultid="648" />
                    <RANKING place="4" resultid="651" />
                    <RANKING place="5" resultid="653" />
                    <RANKING place="1" resultid="663" />
                    <RANKING place="2" resultid="670" />
                    <RANKING place="3" resultid="954" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2" agemax="10" agemin="10" name="Thüringen: Kategorie F (Jg.2013)">
                  <RANKINGS>
                    <RANKING place="1" resultid="266" />
                    <RANKING place="2" resultid="268" />
                    <RANKING place="3" resultid="269" />
                    <RANKING place="5" resultid="270" />
                    <RANKING place="4" resultid="271" />
                    <RANKING place="6" resultid="357" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3" agemax="11" agemin="11" name="Thüringen: Kategorie E (Jg.2012)">
                  <RANKINGS>
                    <RANKING place="1" resultid="264" />
                    <RANKING place="7" resultid="355" />
                    <RANKING place="5" resultid="356" />
                    <RANKING place="8" resultid="362" />
                    <RANKING place="3" resultid="792" />
                    <RANKING place="6" resultid="793" />
                    <RANKING place="2" resultid="794" />
                    <RANKING place="4" resultid="949" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="13" agemin="12" name="Thüringen: Kategorie D (Jg.2010/2011)">
                  <RANKINGS>
                    <RANKING place="3" resultid="263" />
                    <RANKING place="9" resultid="265" />
                    <RANKING place="15" resultid="267" />
                    <RANKING place="2" resultid="359" />
                    <RANKING place="4" resultid="360" />
                    <RANKING place="5" resultid="361" />
                    <RANKING place="10" resultid="607" />
                    <RANKING place="12" resultid="618" />
                    <RANKING place="13" resultid="625" />
                    <RANKING place="16" resultid="780" />
                    <RANKING place="1" resultid="782" />
                    <RANKING place="7" resultid="789" />
                    <RANKING place="17" resultid="791" />
                    <RANKING place="6" resultid="915" />
                    <RANKING place="11" resultid="921" />
                    <RANKING place="8" resultid="927" />
                    <RANKING place="14" resultid="936" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="15" agemin="14" name="Thüringen: Kategorie C (Jg.2008/2009)">
                  <RANKINGS>
                    <RANKING place="6" resultid="511" />
                    <RANKING place="8" resultid="514" />
                    <RANKING place="4" resultid="518" />
                    <RANKING place="3" resultid="596" />
                    <RANKING place="1" resultid="781" />
                    <RANKING place="2" resultid="783" />
                    <RANKING place="5" resultid="902" />
                    <RANKING place="7" resultid="908" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6" agemax="17" agemin="16" name="Thüringen: Kategorie B (Jg.2006/2007)">
                  <RANKINGS>
                    <RANKING place="1" resultid="262" />
                    <RANKING place="3" resultid="491" />
                    <RANKING place="2" resultid="785" />
                    <RANKING place="5" resultid="787" />
                    <RANKING place="4" resultid="888" />
                    <RANKING place="6" resultid="891" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7" agemax="30" agemin="18" name="Thüringen: Kategorie A (Jg.2005 u.ä.)">
                  <RANKINGS>
                    <RANKING place="2" resultid="358" />
                    <RANKING place="1" resultid="565" />
                    <RANKING place="3" resultid="784" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8" agemax="34" agemin="29" name="Thüringen: Master A (Jg.1989-1994)" />
                <AGEGROUP agegroupid="9" agemax="44" agemin="35" name="Thüringen: Master B (Jg.1979-1988)">
                  <RANKINGS>
                    <RANKING place="1" resultid="788" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10" agemax="54" agemin="45" name="Thüringen: Master C (Jg.1969-1978)" />
                <AGEGROUP agegroupid="11" agemax="64" agemin="55" name="Thüringen: Master D (Jg.1959-1968)">
                  <RANKINGS>
                    <RANKING place="1" resultid="790" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="12" agemax="123" agemin="65" name="Thüringen: Master E (Jg.1958 u.ä.)" />
                <AGEGROUP agegroupid="13" agemax="123" agemin="29" name="Offene Wertung Master">
                  <RANKINGS>
                    <RANKING place="3" resultid="677" />
                    <RANKING place="4" resultid="788" />
                    <RANKING place="6" resultid="790" />
                    <RANKING place="2" resultid="825" />
                    <RANKING place="5" resultid="828" />
                    <RANKING place="1" resultid="956" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="14" agemax="30" agemin="1" name="Offene Wertung">
                  <RANKINGS>
                    <RANKING place="3" resultid="32" />
                    <RANKING place="18" resultid="33" />
                    <RANKING place="41" resultid="34" />
                    <RANKING place="46" resultid="35" />
                    <RANKING place="14" resultid="101" />
                    <RANKING place="16" resultid="102" />
                    <RANKING place="23" resultid="103" />
                    <RANKING place="22" resultid="104" />
                    <RANKING place="35" resultid="105" />
                    <RANKING place="29" resultid="106" />
                    <RANKING place="26" resultid="118" />
                    <RANKING place="59" resultid="119" />
                    <RANKING place="2" resultid="129" />
                    <RANKING place="47" resultid="130" />
                    <RANKING place="56" resultid="131" />
                    <RANKING place="64" resultid="132" />
                    <RANKING place="10" resultid="138" />
                    <RANKING place="20" resultid="139" />
                    <RANKING place="4" resultid="180" />
                    <RANKING place="12" resultid="181" />
                    <RANKING place="83" resultid="182" />
                    <RANKING place="89" resultid="183" />
                    <RANKING place="93" resultid="184" />
                    <RANKING place="25" resultid="208" />
                    <RANKING place="8" resultid="262" />
                    <RANKING place="45" resultid="263" />
                    <RANKING place="48" resultid="264" />
                    <RANKING place="61" resultid="265" />
                    <RANKING place="66" resultid="266" />
                    <RANKING place="79" resultid="267" />
                    <RANKING place="82" resultid="268" />
                    <RANKING place="85" resultid="269" />
                    <RANKING place="88" resultid="270" />
                    <RANKING place="86" resultid="271" />
                    <RANKING place="98" resultid="272" />
                    <RANKING place="9" resultid="291" />
                    <RANKING place="75" resultid="292" />
                    <RANKING place="78" resultid="293" />
                    <RANKING place="87" resultid="355" />
                    <RANKING place="76" resultid="356" />
                    <RANKING place="91" resultid="357" />
                    <RANKING place="7" resultid="358" />
                    <RANKING place="42" resultid="359" />
                    <RANKING place="52" resultid="360" />
                    <RANKING place="53" resultid="361" />
                    <RANKING place="90" resultid="362" />
                    <RANKING place="1" resultid="407" />
                    <RANKING place="15" resultid="408" />
                    <RANKING place="12" resultid="456" />
                    <RANKING place="19" resultid="457" />
                    <RANKING place="69" resultid="459" />
                    <RANKING place="74" resultid="460" />
                    <RANKING place="72" resultid="461" />
                    <RANKING place="33" resultid="491" />
                    <RANKING place="49" resultid="511" />
                    <RANKING place="57" resultid="514" />
                    <RANKING place="38" resultid="518" />
                    <RANKING place="36" resultid="537" />
                    <RANKING place="24" resultid="541" />
                    <RANKING place="39" resultid="549" />
                    <RANKING place="44" resultid="553" />
                    <RANKING place="4" resultid="565" />
                    <RANKING place="32" resultid="596" />
                    <RANKING place="63" resultid="607" />
                    <RANKING place="70" resultid="618" />
                    <RANKING place="71" resultid="625" />
                    <RANKING place="99" resultid="648" />
                    <RANKING place="96" resultid="651" />
                    <RANKING place="97" resultid="653" />
                    <RANKING place="92" resultid="663" />
                    <RANKING place="94" resultid="670" />
                    <RANKING place="80" resultid="780" />
                    <RANKING place="11" resultid="781" />
                    <RANKING place="28" resultid="782" />
                    <RANKING place="27" resultid="783" />
                    <RANKING place="37" resultid="784" />
                    <RANKING place="30" resultid="785" />
                    <RANKING place="55" resultid="787" />
                    <RANKING place="58" resultid="789" />
                    <RANKING place="81" resultid="791" />
                    <RANKING place="67" resultid="792" />
                    <RANKING place="84" resultid="793" />
                    <RANKING place="65" resultid="794" />
                    <RANKING place="6" resultid="847" />
                    <RANKING place="17" resultid="850" />
                    <RANKING place="50" resultid="856" />
                    <RANKING place="21" resultid="861" />
                    <RANKING place="31" resultid="865" />
                    <RANKING place="43" resultid="869" />
                    <RANKING place="34" resultid="888" />
                    <RANKING place="62" resultid="891" />
                    <RANKING place="40" resultid="902" />
                    <RANKING place="51" resultid="908" />
                    <RANKING place="54" resultid="915" />
                    <RANKING place="68" resultid="921" />
                    <RANKING place="60" resultid="927" />
                    <RANKING place="77" resultid="936" />
                    <RANKING place="73" resultid="949" />
                    <RANKING place="95" resultid="954" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="12" number="12" gender="M" round="TIM">
              <SWIMSTYLE stroke="SURFACE" relaycount="1" distance="50" />
              <FEE value="500" currency="EUR" />
              <HEATS>
                <HEAT heatid="12001" number="1" />
                <HEAT heatid="12002" number="2" />
                <HEAT heatid="12003" number="3" />
                <HEAT heatid="12004" number="4" />
                <HEAT heatid="12005" number="5" />
                <HEAT heatid="12006" number="6" />
                <HEAT heatid="12007" number="7" />
                <HEAT heatid="12008" number="8" />
                <HEAT heatid="12009" number="9" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="9" agemin="1" name="Thüringen: Kategorie G (Jg.2014 u.j.)">
                  <RANKINGS>
                    <RANKING place="1" resultid="657" />
                    <RANKING place="3" resultid="661" />
                    <RANKING place="4" resultid="666" />
                    <RANKING place="2" resultid="674" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2" agemax="10" agemin="10" name="Thüringen: Kategorie F (Jg.2013)">
                  <RANKINGS>
                    <RANKING place="2" resultid="275" />
                    <RANKING place="3" resultid="364" />
                    <RANKING place="1" resultid="645" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3" agemax="11" agemin="11" name="Thüringen: Kategorie E (Jg.2012)">
                  <RANKINGS>
                    <RANKING place="1" resultid="637" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="13" agemin="12" name="Thüringen: Kategorie D (Jg.2010/2011)">
                  <RANKINGS>
                    <RANKING place="7" resultid="273" />
                    <RANKING place="10" resultid="274" />
                    <RANKING place="1" resultid="369" />
                    <RANKING place="2" resultid="370" />
                    <RANKING place="8" resultid="611" />
                    <RANKING place="4" resultid="799" />
                    <RANKING place="5" resultid="802" />
                    <RANKING place="3" resultid="803" />
                    <RANKING place="6" resultid="805" />
                    <RANKING place="11" resultid="806" />
                    <RANKING place="12" resultid="932" />
                    <RANKING place="9" resultid="941" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="15" agemin="14" name="Thüringen: Kategorie C (Jg.2008/2009)">
                  <RANKINGS>
                    <RANKING place="2" resultid="367" />
                    <RANKING place="7" resultid="373" />
                    <RANKING place="5" resultid="578" />
                    <RANKING place="4" resultid="583" />
                    <RANKING place="1" resultid="587" />
                    <RANKING place="3" resultid="798" />
                    <RANKING place="6" resultid="804" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6" agemax="17" agemin="16" name="Thüringen: Kategorie B (Jg.2006/2007)">
                  <RANKINGS>
                    <RANKING place="2" resultid="366" />
                    <RANKING place="1" resultid="796" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7" agemax="30" agemin="18" name="Thüringen: Kategorie A (Jg.2005 u.ä.)">
                  <RANKINGS>
                    <RANKING place="3" resultid="365" />
                    <RANKING place="1" resultid="880" />
                    <RANKING place="2" resultid="885" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8" agemax="34" agemin="29" name="Thüringen: Master A (Jg.1989-1994)" />
                <AGEGROUP agegroupid="9" agemax="44" agemin="35" name="Thüringen: Master B (Jg.1979-1988)" />
                <AGEGROUP agegroupid="10" agemax="54" agemin="45" name="Thüringen: Master C (Jg.1969-1978)">
                  <RANKINGS>
                    <RANKING place="2" resultid="557" />
                    <RANKING place="1" resultid="797" />
                    <RANKING place="3" resultid="800" />
                    <RANKING place="4" resultid="801" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11" agemax="64" agemin="55" name="Thüringen: Master D (Jg.1959-1968)">
                  <RANKINGS>
                    <RANKING place="1" resultid="371" />
                    <RANKING place="2" resultid="374" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="12" agemax="123" agemin="65" name="Thüringen: Master E (Jg.1958 u.ä.)">
                  <RANKINGS>
                    <RANKING place="1" resultid="372" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="13" agemax="123" agemin="28" name="Offene Wertung Master">
                  <RANKINGS>
                    <RANKING place="5" resultid="371" />
                    <RANKING place="8" resultid="372" />
                    <RANKING place="10" resultid="374" />
                    <RANKING place="4" resultid="557" />
                    <RANKING place="2" resultid="797" />
                    <RANKING place="6" resultid="800" />
                    <RANKING place="9" resultid="801" />
                    <RANKING place="7" resultid="820" />
                    <RANKING place="3" resultid="822" />
                    <RANKING place="1" resultid="958" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="14" agemax="29" agemin="1" name="Offene Wertung">
                  <RANKINGS>
                    <RANKING place="26" resultid="43" />
                    <RANKING place="36" resultid="44" />
                    <RANKING place="1" resultid="51" />
                    <RANKING place="20" resultid="108" />
                    <RANKING place="24" resultid="109" />
                    <RANKING place="29" resultid="110" />
                    <RANKING place="6" resultid="185" />
                    <RANKING place="14" resultid="186" />
                    <RANKING place="53" resultid="187" />
                    <RANKING place="19" resultid="210" />
                    <RANKING place="9" resultid="213" />
                    <RANKING place="41" resultid="273" />
                    <RANKING place="45" resultid="274" />
                    <RANKING place="49" resultid="275" />
                    <RANKING place="57" resultid="364" />
                    <RANKING place="18" resultid="365" />
                    <RANKING place="11" resultid="366" />
                    <RANKING place="16" resultid="367" />
                    <RANKING place="27" resultid="369" />
                    <RANKING place="28" resultid="370" />
                    <RANKING place="37" resultid="373" />
                    <RANKING place="4" resultid="409" />
                    <RANKING place="15" resultid="410" />
                    <RANKING place="22" resultid="412" />
                    <RANKING place="17" resultid="462" />
                    <RANKING place="7" resultid="463" />
                    <RANKING place="21" resultid="464" />
                    <RANKING place="39" resultid="465" />
                    <RANKING place="38" resultid="466" />
                    <RANKING place="42" resultid="467" />
                    <RANKING place="46" resultid="468" />
                    <RANKING place="12" resultid="533" />
                    <RANKING place="25" resultid="545" />
                    <RANKING place="34" resultid="578" />
                    <RANKING place="33" resultid="583" />
                    <RANKING place="10" resultid="587" />
                    <RANKING place="43" resultid="611" />
                    <RANKING place="47" resultid="637" />
                    <RANKING place="48" resultid="645" />
                    <RANKING place="51" resultid="657" />
                    <RANKING place="55" resultid="661" />
                    <RANKING place="56" resultid="666" />
                    <RANKING place="54" resultid="674" />
                    <RANKING place="2" resultid="796" />
                    <RANKING place="23" resultid="798" />
                    <RANKING place="31" resultid="799" />
                    <RANKING place="32" resultid="802" />
                    <RANKING place="30" resultid="803" />
                    <RANKING place="35" resultid="804" />
                    <RANKING place="40" resultid="805" />
                    <RANKING place="50" resultid="806" />
                    <RANKING place="5" resultid="834" />
                    <RANKING place="8" resultid="842" />
                    <RANKING place="3" resultid="880" />
                    <RANKING place="13" resultid="885" />
                    <RANKING place="52" resultid="932" />
                    <RANKING place="44" resultid="941" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="13" number="13" gender="F" round="TIM">
              <SWIMSTYLE stroke="SURFACE" relaycount="1" distance="200" />
              <FEE value="500" currency="EUR" />
              <HEATS>
                <HEAT heatid="13001" number="1" />
                <HEAT heatid="13002" number="2" />
                <HEAT heatid="13003" number="3" />
                <HEAT heatid="13004" number="4" />
                <HEAT heatid="13005" number="5" />
                <HEAT heatid="13006" number="6" />
                <HEAT heatid="13007" number="7" />
                <HEAT heatid="13008" number="8" />
                <HEAT heatid="13009" number="9" />
                <HEAT heatid="13010" number="10" />
                <HEAT heatid="13011" number="11" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="9" agemin="1" name="Thüringen: Kategorie G (Jg.2014 u.j.)">
                  <RANKINGS>
                    <RANKING place="1" resultid="526" />
                    <RANKING place="3" resultid="649" />
                    <RANKING place="2" resultid="961" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2" agemax="10" agemin="10" name="Thüringen: Kategorie F (Jg.2013)">
                  <RANKINGS>
                    <RANKING place="3" resultid="236" />
                    <RANKING place="2" resultid="241" />
                    <RANKING place="1" resultid="242" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3" agemax="11" agemin="11" name="Thüringen: Kategorie E (Jg.2012)">
                  <RANKINGS>
                    <RANKING place="1" resultid="240" />
                    <RANKING place="2" resultid="737" />
                    <RANKING place="3" resultid="738" />
                    <RANKING place="4" resultid="950" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="13" agemin="12" name="Thüringen: Kategorie D (Jg.2010/2011)">
                  <RANKINGS>
                    <RANKING place="7" resultid="233" />
                    <RANKING place="14" resultid="235" />
                    <RANKING place="2" resultid="239" />
                    <RANKING place="6" resultid="321" />
                    <RANKING place="13" resultid="322" />
                    <RANKING place="3" resultid="323" />
                    <RANKING place="10" resultid="608" />
                    <RANKING place="9" resultid="619" />
                    <RANKING place="11" resultid="626" />
                    <RANKING place="15" resultid="729" />
                    <RANKING place="1" resultid="731" />
                    <RANKING place="8" resultid="736" />
                    <RANKING place="4" resultid="916" />
                    <RANKING place="12" resultid="922" />
                    <RANKING place="5" resultid="928" />
                    <RANKING place="16" resultid="937" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="15" agemin="14" name="Thüringen: Kategorie C (Jg.2008/2009)">
                  <RANKINGS>
                    <RANKING place="4" resultid="507" />
                    <RANKING place="5" resultid="515" />
                    <RANKING place="2" resultid="591" />
                    <RANKING place="1" resultid="732" />
                    <RANKING place="3" resultid="909" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6" agemax="17" agemin="16" name="Thüringen: Kategorie B (Jg.2006/2007)">
                  <RANKINGS>
                    <RANKING place="3" resultid="238" />
                    <RANKING place="2" resultid="492" />
                    <RANKING place="1" resultid="733" />
                    <RANKING place="4" resultid="735" />
                    <RANKING place="5" resultid="892" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7" agemax="30" agemin="18" name="Thüringen: Kategorie A (Jg.2005 u.ä.)">
                  <RANKINGS>
                    <RANKING place="2" resultid="237" />
                    <RANKING place="1" resultid="566" />
                    <RANKING place="3" resultid="730" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8" agemax="34" agemin="29" name="Thüringen: Master A (Jg.1989-1994)" />
                <AGEGROUP agegroupid="9" agemax="44" agemin="35" name="Thüringen: Master B (Jg.1979-1988)" />
                <AGEGROUP agegroupid="10" agemax="54" agemin="45" name="Thüringen: Master C (Jg.1969-1978)" />
                <AGEGROUP agegroupid="11" agemax="64" agemin="55" name="Thüringen: Master D (Jg.1959-1968)" />
                <AGEGROUP agegroupid="12" agemax="123" agemin="65" name="Thüringen: Master E (Jg.1958 u.ä.)" />
                <AGEGROUP agegroupid="13" agemax="123" agemin="29" name="Offene Wertung Master">
                  <RANKINGS>
                    <RANKING place="1" resultid="826" />
                    <RANKING place="2" resultid="829" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="14" agemax="30" agemin="1" name="Offene Wertung">
                  <RANKINGS>
                    <RANKING place="5" resultid="10" />
                    <RANKING place="9" resultid="11" />
                    <RANKING place="39" resultid="12" />
                    <RANKING place="36" resultid="13" />
                    <RANKING place="19" resultid="74" />
                    <RANKING place="13" resultid="75" />
                    <RANKING place="24" resultid="76" />
                    <RANKING place="34" resultid="77" />
                    <RANKING place="32" resultid="78" />
                    <RANKING place="41" resultid="79" />
                    <RANKING place="51" resultid="115" />
                    <RANKING place="2" resultid="154" />
                    <RANKING place="3" resultid="155" />
                    <RANKING place="14" resultid="156" />
                    <RANKING place="6" resultid="157" />
                    <RANKING place="17" resultid="158" />
                    <RANKING place="18" resultid="159" />
                    <RANKING place="15" resultid="214" />
                    <RANKING place="52" resultid="233" />
                    <RANKING place="71" resultid="235" />
                    <RANKING place="72" resultid="236" />
                    <RANKING place="16" resultid="237" />
                    <RANKING place="33" resultid="238" />
                    <RANKING place="46" resultid="239" />
                    <RANKING place="43" resultid="240" />
                    <RANKING place="66" resultid="241" />
                    <RANKING place="61" resultid="242" />
                    <RANKING place="8" resultid="283" />
                    <RANKING place="65" resultid="284" />
                    <RANKING place="69" resultid="285" />
                    <RANKING place="50" resultid="321" />
                    <RANKING place="60" resultid="322" />
                    <RANKING place="47" resultid="323" />
                    <RANKING place="4" resultid="390" />
                    <RANKING place="12" resultid="391" />
                    <RANKING place="10" resultid="425" />
                    <RANKING place="20" resultid="426" />
                    <RANKING place="27" resultid="427" />
                    <RANKING place="28" resultid="428" />
                    <RANKING place="67" resultid="429" />
                    <RANKING place="70" resultid="430" />
                    <RANKING place="68" resultid="431" />
                    <RANKING place="75" resultid="432" />
                    <RANKING place="31" resultid="492" />
                    <RANKING place="45" resultid="507" />
                    <RANKING place="55" resultid="515" />
                    <RANKING place="76" resultid="526" />
                    <RANKING place="11" resultid="566" />
                    <RANKING place="37" resultid="591" />
                    <RANKING place="57" resultid="608" />
                    <RANKING place="56" resultid="619" />
                    <RANKING place="58" resultid="626" />
                    <RANKING place="78" resultid="649" />
                    <RANKING place="1" resultid="681" />
                    <RANKING place="7" resultid="685" />
                    <RANKING place="23" resultid="688" />
                    <RANKING place="73" resultid="729" />
                    <RANKING place="22" resultid="730" />
                    <RANKING place="25" resultid="731" />
                    <RANKING place="30" resultid="732" />
                    <RANKING place="26" resultid="733" />
                    <RANKING place="44" resultid="735" />
                    <RANKING place="53" resultid="736" />
                    <RANKING place="54" resultid="737" />
                    <RANKING place="63" resultid="738" />
                    <RANKING place="21" resultid="851" />
                    <RANKING place="38" resultid="857" />
                    <RANKING place="29" resultid="862" />
                    <RANKING place="35" resultid="866" />
                    <RANKING place="40" resultid="870" />
                    <RANKING place="62" resultid="892" />
                    <RANKING place="42" resultid="909" />
                    <RANKING place="48" resultid="916" />
                    <RANKING place="59" resultid="922" />
                    <RANKING place="49" resultid="928" />
                    <RANKING place="74" resultid="937" />
                    <RANKING place="64" resultid="950" />
                    <RANKING place="77" resultid="961" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="14" number="14" gender="M" round="TIM">
              <SWIMSTYLE stroke="SURFACE" relaycount="1" distance="200" />
              <FEE value="500" currency="EUR" />
              <HEATS>
                <HEAT heatid="14001" number="1" />
                <HEAT heatid="14002" number="2" />
                <HEAT heatid="14003" number="3" />
                <HEAT heatid="14004" number="4" />
                <HEAT heatid="14005" number="5" />
                <HEAT heatid="14006" number="6" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="9" agemin="1" name="Thüringen: Kategorie G (Jg.2014 u.j.)">
                  <RANKINGS>
                    <RANKING place="1" resultid="667" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2" agemax="10" agemin="10" name="Thüringen: Kategorie F (Jg.2013)">
                  <RANKINGS>
                    <RANKING place="2" resultid="243" />
                    <RANKING place="1" resultid="646" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3" agemax="11" agemin="11" name="Thüringen: Kategorie E (Jg.2012)">
                  <RANKINGS>
                    <RANKING place="2" resultid="521" />
                    <RANKING place="1" resultid="638" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="13" agemin="12" name="Thüringen: Kategorie D (Jg.2010/2011)">
                  <RANKINGS>
                    <RANKING place="8" resultid="244" />
                    <RANKING place="7" resultid="245" />
                    <RANKING place="6" resultid="325" />
                    <RANKING place="2" resultid="327" />
                    <RANKING place="5" resultid="622" />
                    <RANKING place="1" resultid="740" />
                    <RANKING place="4" resultid="741" />
                    <RANKING place="3" resultid="742" />
                    <RANKING place="9" resultid="745" />
                    <RANKING place="11" resultid="933" />
                    <RANKING place="10" resultid="942" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="15" agemin="14" name="Thüringen: Kategorie C (Jg.2008/2009)">
                  <RANKINGS>
                    <RANKING place="7" resultid="326" />
                    <RANKING place="2" resultid="502" />
                    <RANKING place="5" resultid="584" />
                    <RANKING place="1" resultid="588" />
                    <RANKING place="3" resultid="601" />
                    <RANKING place="4" resultid="739" />
                    <RANKING place="6" resultid="743" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6" agemax="17" agemin="16" name="Thüringen: Kategorie B (Jg.2006/2007)">
                  <RANKINGS>
                    <RANKING place="1" resultid="500" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7" agemax="30" agemin="18" name="Thüringen: Kategorie A (Jg.2005 u.ä.)">
                  <RANKINGS>
                    <RANKING place="1" resultid="324" />
                    <RANKING place="2" resultid="881" />
                    <RANKING place="3" resultid="886" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8" agemax="34" agemin="29" name="Thüringen: Master A (Jg.1989-1994)" />
                <AGEGROUP agegroupid="9" agemax="44" agemin="35" name="Thüringen: Master B (Jg.1979-1988)" />
                <AGEGROUP agegroupid="10" agemax="54" agemin="45" name="Thüringen: Master C (Jg.1969-1978)" />
                <AGEGROUP agegroupid="11" agemax="64" agemin="55" name="Thüringen: Master D (Jg.1959-1968)" />
                <AGEGROUP agegroupid="12" agemax="123" agemin="65" name="Thüringen: Master E (Jg.1958 u.ä.)" />
                <AGEGROUP agegroupid="13" agemax="123" agemin="28" name="Offene Wertung Master">
                  <RANKINGS>
                    <RANKING place="1" resultid="959" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="14" agemax="29" agemin="1" name="Offene Wertung">
                  <RANKINGS>
                    <RANKING place="2" resultid="14" />
                    <RANKING place="5" resultid="15" />
                    <RANKING place="14" resultid="16" />
                    <RANKING place="20" resultid="38" />
                    <RANKING place="10" resultid="80" />
                    <RANKING place="12" resultid="81" />
                    <RANKING place="19" resultid="82" />
                    <RANKING place="3" resultid="160" />
                    <RANKING place="11" resultid="162" />
                    <RANKING place="40" resultid="243" />
                    <RANKING place="34" resultid="244" />
                    <RANKING place="32" resultid="245" />
                    <RANKING place="4" resultid="324" />
                    <RANKING place="31" resultid="325" />
                    <RANKING place="26" resultid="326" />
                    <RANKING place="21" resultid="327" />
                    <RANKING place="1" resultid="392" />
                    <RANKING place="13" resultid="433" />
                    <RANKING place="30" resultid="434" />
                    <RANKING place="29" resultid="436" />
                    <RANKING place="27" resultid="500" />
                    <RANKING place="15" resultid="502" />
                    <RANKING place="37" resultid="521" />
                    <RANKING place="22" resultid="584" />
                    <RANKING place="8" resultid="588" />
                    <RANKING place="16" resultid="601" />
                    <RANKING place="28" resultid="622" />
                    <RANKING place="33" resultid="638" />
                    <RANKING place="35" resultid="646" />
                    <RANKING place="41" resultid="667" />
                    <RANKING place="18" resultid="739" />
                    <RANKING place="17" resultid="740" />
                    <RANKING place="25" resultid="741" />
                    <RANKING place="24" resultid="742" />
                    <RANKING place="23" resultid="743" />
                    <RANKING place="36" resultid="745" />
                    <RANKING place="6" resultid="835" />
                    <RANKING place="7" resultid="881" />
                    <RANKING place="9" resultid="886" />
                    <RANKING place="39" resultid="933" />
                    <RANKING place="38" resultid="942" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="15" number="15" gender="X" round="TIM">
              <SWIMSTYLE stroke="SURFACE" relaycount="4" distance="50" />
              <FEE value="800" currency="EUR" />
              <HEATS>
                <HEAT heatid="15001" number="1" />
                <HEAT heatid="15002" number="2" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="11" agemin="1" name="Thüringen: Kategorie III (Jg.2012 u.j.)">
                  <RANKINGS>
                    <RANKING place="1" resultid="255" />
                    <RANKING place="3" resultid="256" />
                    <RANKING place="5" resultid="336" />
                    <RANKING place="4" resultid="634" />
                    <RANKING place="7" resultid="654" />
                    <RANKING place="6" resultid="671" />
                    <RANKING place="2" resultid="763" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="11" agemin="1" name="Offene Wertung">
                  <RANKINGS>
                    <RANKING place="6" resultid="170" />
                    <RANKING place="1" resultid="255" />
                    <RANKING place="3" resultid="256" />
                    <RANKING place="5" resultid="336" />
                    <RANKING place="4" resultid="634" />
                    <RANKING place="8" resultid="654" />
                    <RANKING place="7" resultid="671" />
                    <RANKING place="2" resultid="763" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2" agemax="-1" agemin="180" easy.ak="180" calculate="TOTAL" name="Thüringen: Master I (Gesamtalter &lt;= 180 Jahre)">
                  <RANKINGS>
                    <RANKING place="1" resultid="762" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3" agemax="-1" agemin="400" easy.ak="400" calculate="TOTAL" name="Thüringen: Master II (Gesamtalter &gt; 181 Jahre)">
                  <RANKINGS>
                    <RANKING place="1" resultid="337" />
                    <RANKING place="2" resultid="761" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="-1" agemin="400" easy.ak="400" calculate="TOTAL" name="Offene Wertung Master">
                  <RANKINGS>
                    <RANKING place="1" resultid="337" />
                    <RANKING place="3" resultid="761" />
                    <RANKING place="4" resultid="762" />
                    <RANKING place="2" resultid="817" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="16" number="16" gender="F" round="TIM">
              <SWIMSTYLE stroke="SURFACE" relaycount="1" distance="400" />
              <FEE value="500" currency="EUR" />
              <HEATS>
                <HEAT heatid="16001" number="1" />
                <HEAT heatid="16002" number="2" />
                <HEAT heatid="16003" number="3" />
                <HEAT heatid="16004" number="4" />
                <HEAT heatid="16005" number="5" />
                <HEAT heatid="16006" number="6" />
                <HEAT heatid="16007" number="7" />
                <HEAT heatid="16008" number="8" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="9" agemin="10" name="Thüringen: Kategorie G (Jg.2014 u.j.)" />
                <AGEGROUP agegroupid="2" agemax="10" agemin="10" name="Thüringen: Kategorie F (Jg.2013)">
                  <RANKINGS>
                    <RANKING place="2" resultid="246" />
                    <RANKING place="1" resultid="247" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3" agemax="11" agemin="11" name="Thüringen: Kategorie E (Jg.2012)">
                  <RANKINGS>
                    <RANKING place="1" resultid="249" />
                    <RANKING place="2" resultid="749" />
                    <RANKING place="3" resultid="951" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="13" agemin="12" name="Thüringen: Kategorie D (Jg.2010/2011)">
                  <RANKINGS>
                    <RANKING place="1" resultid="329" />
                    <RANKING place="4" resultid="627" />
                    <RANKING place="7" resultid="750" />
                    <RANKING place="3" resultid="917" />
                    <RANKING place="5" resultid="923" />
                    <RANKING place="2" resultid="929" />
                    <RANKING place="6" resultid="938" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="15" agemin="14" name="Thüringen: Kategorie C (Jg.2008/2009)">
                  <RANKINGS>
                    <RANKING place="3" resultid="512" />
                    <RANKING place="4" resultid="519" />
                    <RANKING place="1" resultid="748" />
                    <RANKING place="2" resultid="903" />
                    <RANKING place="5" resultid="910" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6" agemax="17" agemin="16" name="Thüringen: Kategorie B (Jg.2006/2007)">
                  <RANKINGS>
                    <RANKING place="1" resultid="893" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7" agemax="30" agemin="18" name="Thüringen: Kategorie A (Jg.2005 u.ä.)">
                  <RANKINGS>
                    <RANKING place="2" resultid="330" />
                    <RANKING place="4" resultid="476" />
                    <RANKING place="1" resultid="480" />
                    <RANKING place="3" resultid="567" />
                    <RANKING place="5" resultid="747" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8" agemax="34" agemin="29" name="Thüringen: Master A (Jg.1989-1994)" />
                <AGEGROUP agegroupid="9" agemax="44" agemin="35" name="Thüringen: Master B (Jg.1979-1988)" />
                <AGEGROUP agegroupid="10" agemax="54" agemin="45" name="Thüringen: Master C (Jg.1969-1978)" />
                <AGEGROUP agegroupid="11" agemax="64" agemin="55" name="Thüringen: Master D (Jg.1959-1968)" />
                <AGEGROUP agegroupid="12" agemax="123" agemin="65" name="Thüringen: Master E (Jg.1958 u.ä.)" />
                <AGEGROUP agegroupid="13" agemax="123" agemin="29" name="Offene Wertung Master">
                  <RANKINGS>
                    <RANKING place="1" resultid="830" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="14" agemax="30" agemin="10" name="Offene Wertung">
                  <RANKINGS>
                    <RANKING place="4" resultid="17" />
                    <RANKING place="8" resultid="18" />
                    <RANKING place="16" resultid="54" />
                    <RANKING place="24" resultid="83" />
                    <RANKING place="28" resultid="84" />
                    <RANKING place="29" resultid="85" />
                    <RANKING place="41" resultid="86" />
                    <RANKING place="12" resultid="126" />
                    <RANKING place="34" resultid="136" />
                    <RANKING place="2" resultid="163" />
                    <RANKING place="14" resultid="164" />
                    <RANKING place="9" resultid="165" />
                    <RANKING place="20" resultid="166" />
                    <RANKING place="27" resultid="200" />
                    <RANKING place="54" resultid="246" />
                    <RANKING place="51" resultid="247" />
                    <RANKING place="43" resultid="249" />
                    <RANKING place="7" resultid="286" />
                    <RANKING place="3" resultid="287" />
                    <RANKING place="44" resultid="329" />
                    <RANKING place="13" resultid="330" />
                    <RANKING place="1" resultid="393" />
                    <RANKING place="6" resultid="394" />
                    <RANKING place="10" resultid="395" />
                    <RANKING place="19" resultid="396" />
                    <RANKING place="21" resultid="438" />
                    <RANKING place="17" resultid="439" />
                    <RANKING place="26" resultid="440" />
                    <RANKING place="18" resultid="476" />
                    <RANKING place="11" resultid="480" />
                    <RANKING place="35" resultid="512" />
                    <RANKING place="38" resultid="519" />
                    <RANKING place="32" resultid="542" />
                    <RANKING place="39" resultid="550" />
                    <RANKING place="37" resultid="554" />
                    <RANKING place="15" resultid="567" />
                    <RANKING place="48" resultid="627" />
                    <RANKING place="22" resultid="689" />
                    <RANKING place="23" resultid="747" />
                    <RANKING place="30" resultid="748" />
                    <RANKING place="47" resultid="749" />
                    <RANKING place="55" resultid="750" />
                    <RANKING place="5" resultid="848" />
                    <RANKING place="36" resultid="858" />
                    <RANKING place="25" resultid="863" />
                    <RANKING place="31" resultid="867" />
                    <RANKING place="40" resultid="871" />
                    <RANKING place="50" resultid="893" />
                    <RANKING place="33" resultid="903" />
                    <RANKING place="42" resultid="910" />
                    <RANKING place="46" resultid="917" />
                    <RANKING place="49" resultid="923" />
                    <RANKING place="45" resultid="929" />
                    <RANKING place="53" resultid="938" />
                    <RANKING place="52" resultid="951" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="17" number="17" gender="M" round="TIM">
              <SWIMSTYLE stroke="SURFACE" relaycount="1" distance="400" />
              <FEE value="500" currency="EUR" />
              <HEATS>
                <HEAT heatid="17001" number="1" />
                <HEAT heatid="17002" number="2" />
                <HEAT heatid="17003" number="3" />
                <HEAT heatid="17004" number="4" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="9" agemin="10" name="Thüringen: Kategorie G (Jg.2014 u.j.)" />
                <AGEGROUP agegroupid="2" agemax="10" agemin="10" name="Thüringen: Kategorie F (Jg.2013)" />
                <AGEGROUP agegroupid="3" agemax="11" agemin="11" name="Thüringen: Kategorie E (Jg.2012)">
                  <RANKINGS>
                    <RANKING place="2" resultid="522" />
                    <RANKING place="1" resultid="639" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="13" agemin="12" name="Thüringen: Kategorie D (Jg.2010/2011)">
                  <RANKINGS>
                    <RANKING place="4" resultid="250" />
                    <RANKING place="2" resultid="623" />
                    <RANKING place="1" resultid="752" />
                    <RANKING place="3" resultid="753" />
                    <RANKING place="6" resultid="934" />
                    <RANKING place="5" resultid="943" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="15" agemin="14" name="Thüringen: Kategorie C (Jg.2008/2009)">
                  <RANKINGS>
                    <RANKING place="1" resultid="503" />
                    <RANKING place="2" resultid="602" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6" agemax="17" agemin="16" name="Thüringen: Kategorie B (Jg.2006/2007)">
                  <RANKINGS>
                    <RANKING place="1" resultid="898" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7" agemax="30" agemin="18" name="Thüringen: Kategorie A (Jg.2005 u.ä.)" />
                <AGEGROUP agegroupid="8" agemax="34" agemin="29" name="Thüringen: Master A (Jg.1989-1994)" />
                <AGEGROUP agegroupid="9" agemax="44" agemin="35" name="Thüringen: Master B (Jg.1979-1988)" />
                <AGEGROUP agegroupid="10" agemax="54" agemin="45" name="Thüringen: Master C (Jg.1969-1978)" />
                <AGEGROUP agegroupid="11" agemax="64" agemin="55" name="Thüringen: Master D (Jg.1959-1968)" />
                <AGEGROUP agegroupid="12" agemax="123" agemin="65" name="Thüringen: Master E (Jg.1958 u.ä.)" />
                <AGEGROUP agegroupid="13" agemax="123" agemin="28" name="Offene Wertung Master">
                  <RANKINGS>
                    <RANKING place="1" resultid="960" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="14" agemax="29" agemin="10" name="Offene Wertung">
                  <RANKINGS>
                    <RANKING place="5" resultid="20" />
                    <RANKING place="7" resultid="21" />
                    <RANKING place="13" resultid="39" />
                    <RANKING place="16" resultid="40" />
                    <RANKING place="4" resultid="49" />
                    <RANKING place="11" resultid="87" />
                    <RANKING place="9" resultid="88" />
                    <RANKING place="21" resultid="250" />
                    <RANKING place="1" resultid="398" />
                    <RANKING place="3" resultid="399" />
                    <RANKING place="6" resultid="401" />
                    <RANKING place="8" resultid="441" />
                    <RANKING place="10" resultid="503" />
                    <RANKING place="22" resultid="522" />
                    <RANKING place="2" resultid="529" />
                    <RANKING place="12" resultid="546" />
                    <RANKING place="14" resultid="602" />
                    <RANKING place="18" resultid="623" />
                    <RANKING place="20" resultid="639" />
                    <RANKING place="17" resultid="752" />
                    <RANKING place="19" resultid="753" />
                    <RANKING place="15" resultid="898" />
                    <RANKING place="24" resultid="934" />
                    <RANKING place="23" resultid="943" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="18" number="18" gender="F" round="TIM">
              <SWIMSTYLE stroke="IMMERSION" technique="DIVE" relaycount="1" distance="100" />
              <FEE value="500" currency="EUR" />
              <HEATS>
                <HEAT heatid="18001" number="1" />
                <HEAT heatid="18002" number="2" />
                <HEAT heatid="18003" number="3" />
                <HEAT heatid="18004" number="4" />
                <HEAT heatid="18005" number="5" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="9" agemin="12" name="Thüringen: Kategorie G (Jg.2014 u.j.)" />
                <AGEGROUP agegroupid="2" agemax="10" agemin="12" name="Thüringen: Kategorie F (Jg.2013)" />
                <AGEGROUP agegroupid="3" agemax="11" agemin="12" name="Thüringen: Kategorie E (Jg.2012)" />
                <AGEGROUP agegroupid="4" agemax="13" agemin="12" name="Thüringen: Kategorie D (Jg.2010/2011)">
                  <RANKINGS>
                    <RANKING place="2" resultid="230" />
                    <RANKING place="1" resultid="720" />
                    <RANKING place="3" resultid="918" />
                    <RANKING place="4" resultid="924" />
                    <RANKING place="5" resultid="930" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="15" agemin="14" name="Thüringen: Kategorie C (Jg.2008/2009)">
                  <RANKINGS>
                    <RANKING place="6" resultid="508" />
                    <RANKING place="7" resultid="516" />
                    <RANKING place="3" resultid="520" />
                    <RANKING place="1" resultid="592" />
                    <RANKING place="2" resultid="721" />
                    <RANKING place="4" resultid="904" />
                    <RANKING place="5" resultid="911" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6" agemax="17" agemin="16" name="Thüringen: Kategorie B (Jg.2006/2007)">
                  <RANKINGS>
                    <RANKING place="2" resultid="232" />
                    <RANKING place="4" resultid="493" />
                    <RANKING place="5" resultid="496" />
                    <RANKING place="1" resultid="572" />
                    <RANKING place="3" resultid="722" />
                    <RANKING place="6" resultid="894" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7" agemax="30" agemin="18" name="Thüringen: Kategorie A (Jg.2005 u.ä.)">
                  <RANKINGS>
                    <RANKING place="2" resultid="231" />
                    <RANKING place="1" resultid="314" />
                    <RANKING place="3" resultid="481" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8" agemax="34" agemin="29" name="Thüringen: Master A (Jg.1989-1994)" />
                <AGEGROUP agegroupid="9" agemax="44" agemin="35" name="Thüringen: Master B (Jg.1979-1988)" />
                <AGEGROUP agegroupid="10" agemax="54" agemin="45" name="Thüringen: Master C (Jg.1969-1978)" />
                <AGEGROUP agegroupid="11" agemax="64" agemin="55" name="Thüringen: Master D (Jg.1959-1968)" />
                <AGEGROUP agegroupid="12" agemax="123" agemin="65" name="Thüringen: Master E (Jg.1958 u.ä.)" />
                <AGEGROUP agegroupid="13" agemax="123" agemin="29" name="Offene Wertung Master">
                  <RANKINGS>
                    <RANKING place="1" resultid="678" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="14" agemax="30" agemin="12" name="Offene Wertung">
                  <RANKINGS>
                    <RANKING place="11" resultid="53" />
                    <RANKING place="15" resultid="69" />
                    <RANKING place="17" resultid="70" />
                    <RANKING place="21" resultid="114" />
                    <RANKING place="3" resultid="124" />
                    <RANKING place="33" resultid="125" />
                    <RANKING place="5" resultid="135" />
                    <RANKING place="9" resultid="150" />
                    <RANKING place="12" resultid="195" />
                    <RANKING place="14" resultid="196" />
                    <RANKING place="30" resultid="230" />
                    <RANKING place="6" resultid="231" />
                    <RANKING place="13" resultid="232" />
                    <RANKING place="4" resultid="314" />
                    <RANKING place="10" resultid="387" />
                    <RANKING place="16" resultid="388" />
                    <RANKING place="7" resultid="481" />
                    <RANKING place="25" resultid="493" />
                    <RANKING place="28" resultid="496" />
                    <RANKING place="31" resultid="508" />
                    <RANKING place="37" resultid="516" />
                    <RANKING place="26" resultid="520" />
                    <RANKING place="24" resultid="538" />
                    <RANKING place="8" resultid="572" />
                    <RANKING place="20" resultid="592" />
                    <RANKING place="1" resultid="682" />
                    <RANKING place="2" resultid="686" />
                    <RANKING place="23" resultid="720" />
                    <RANKING place="22" resultid="721" />
                    <RANKING place="19" resultid="722" />
                    <RANKING place="18" resultid="852" />
                    <RANKING place="34" resultid="894" />
                    <RANKING place="27" resultid="904" />
                    <RANKING place="29" resultid="911" />
                    <RANKING place="32" resultid="918" />
                    <RANKING place="35" resultid="924" />
                    <RANKING place="36" resultid="930" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="19" number="19" gender="M" round="TIM">
              <SWIMSTYLE stroke="IMMERSION" technique="DIVE" relaycount="1" distance="100" />
              <FEE value="500" currency="EUR" />
              <HEATS>
                <HEAT heatid="19001" number="1" />
                <HEAT heatid="19002" number="2" />
                <HEAT heatid="19003" number="3" />
                <HEAT heatid="19004" number="4" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="9" agemin="12" name="Thüringen: Kategorie G (Jg.2014 u.j.)" />
                <AGEGROUP agegroupid="2" agemax="10" agemin="12" name="Thüringen: Kategorie F (Jg.2013)" />
                <AGEGROUP agegroupid="3" agemax="11" agemin="12" name="Thüringen: Kategorie E (Jg.2012)" />
                <AGEGROUP agegroupid="4" agemax="13" agemin="12" name="Thüringen: Kategorie D (Jg.2010/2011)">
                  <RANKINGS>
                    <RANKING place="2" resultid="319" />
                    <RANKING place="3" resultid="320" />
                    <RANKING place="1" resultid="726" />
                    <RANKING place="4" resultid="944" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="15" agemin="14" name="Thüringen: Kategorie C (Jg.2008/2009)">
                  <RANKINGS>
                    <RANKING place="1" resultid="317" />
                    <RANKING place="3" resultid="504" />
                    <RANKING place="7" resultid="580" />
                    <RANKING place="6" resultid="585" />
                    <RANKING place="2" resultid="589" />
                    <RANKING place="5" resultid="603" />
                    <RANKING place="8" resultid="723" />
                    <RANKING place="4" resultid="727" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6" agemax="17" agemin="16" name="Thüringen: Kategorie B (Jg.2006/2007)">
                  <RANKINGS>
                    <RANKING place="1" resultid="724" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7" agemax="44" agemin="18" name="Thüringen: Kategorie A (Jg.2005 u.ä.)">
                  <RANKINGS>
                    <RANKING place="1" resultid="315" />
                    <RANKING place="3" resultid="316" />
                    <RANKING place="4" resultid="472" />
                    <RANKING place="2" resultid="877" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8" agemax="34" agemin="29" name="Thüringen: Master A (Jg.1989-1994)" />
                <AGEGROUP agegroupid="9" agemax="43" agemin="35" name="Thüringen: Master B (Jg.1979-1988)" />
                <AGEGROUP agegroupid="10" agemax="54" agemin="45" name="Thüringen: Master C (Jg.1969-1978)">
                  <RANKINGS>
                    <RANKING place="1" resultid="725" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11" agemax="64" agemin="55" name="Thüringen: Master D (Jg.1959-1968)" />
                <AGEGROUP agegroupid="12" agemax="123" agemin="65" name="Thüringen: Master E (Jg.1958 u.ä.)" />
                <AGEGROUP agegroupid="13" agemax="123" agemin="45" name="Offene Wertung Master">
                  <RANKINGS>
                    <RANKING place="1" resultid="725" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="14" agemax="44" agemin="12" name="Offene Wertung">
                  <RANKINGS>
                    <RANKING place="3" resultid="9" />
                    <RANKING place="13" resultid="72" />
                    <RANKING place="17" resultid="73" />
                    <RANKING place="7" resultid="151" />
                    <RANKING place="2" resultid="197" />
                    <RANKING place="4" resultid="315" />
                    <RANKING place="12" resultid="316" />
                    <RANKING place="6" resultid="317" />
                    <RANKING place="19" resultid="319" />
                    <RANKING place="22" resultid="320" />
                    <RANKING place="24" resultid="472" />
                    <RANKING place="14" resultid="504" />
                    <RANKING place="5" resultid="530" />
                    <RANKING place="10" resultid="534" />
                    <RANKING place="21" resultid="580" />
                    <RANKING place="20" resultid="585" />
                    <RANKING place="9" resultid="589" />
                    <RANKING place="16" resultid="603" />
                    <RANKING place="23" resultid="723" />
                    <RANKING place="1" resultid="724" />
                    <RANKING place="18" resultid="726" />
                    <RANKING place="15" resultid="727" />
                    <RANKING place="11" resultid="843" />
                    <RANKING place="8" resultid="877" />
                    <RANKING place="25" resultid="944" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="20" number="20" gender="F" round="TIM">
              <SWIMSTYLE stroke="SURFACE" relaycount="4" distance="100" />
              <FEE value="800" currency="EUR" />
              <HEATS>
                <HEAT heatid="20001" number="1" />
                <HEAT heatid="20002" number="2" />
                <HEAT heatid="20003" number="3" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="11" agemin="1" name="Thüringen: Kategorie III (Jg.2012 u.j.)">
                  <RANKINGS>
                    <RANKING place="1" resultid="252" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2" agemax="17" agemin="12" name="Thüringen: Kategorie II (Jg.2006-2011)">
                  <RANKINGS>
                    <RANKING place="5" resultid="253" />
                    <RANKING place="2" resultid="497" />
                    <RANKING place="1" resultid="754" />
                    <RANKING place="4" resultid="756" />
                    <RANKING place="3" resultid="912" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3" agemax="123" agemin="18" name="Thüringen: Kategorie I (Jg.2005 u.ä.)">
                  <RANKINGS>
                    <RANKING place="1" resultid="477" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="123" agemin="1" name="Offene Wertung">
                  <RANKINGS>
                    <RANKING place="2" resultid="23" />
                    <RANKING place="7" resultid="89" />
                    <RANKING place="5" resultid="127" />
                    <RANKING place="13" resultid="252" />
                    <RANKING place="15" resultid="253" />
                    <RANKING place="10" resultid="288" />
                    <RANKING place="1" resultid="402" />
                    <RANKING place="3" resultid="442" />
                    <RANKING place="14" resultid="443" />
                    <RANKING place="6" resultid="477" />
                    <RANKING place="9" resultid="497" />
                    <RANKING place="4" resultid="754" />
                    <RANKING place="12" resultid="756" />
                    <RANKING place="8" resultid="853" />
                    <RANKING place="11" resultid="912" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="21" number="21" gender="X" round="TIM">
              <SWIMSTYLE stroke="SURFACE" relaycount="4" distance="100" />
              <FEE value="800" currency="EUR" />
              <HEATS>
                <HEAT heatid="21001" number="1" />
                <HEAT heatid="21002" number="2" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="5" agemax="11" agemin="1" name="Thüringen: Kategorie III (Jg.2012 u.j.)" />
                <AGEGROUP agegroupid="6" agemax="17" agemin="12" name="Thüringen: Kategorie II (Jg.2006-2011)">
                  <RANKINGS>
                    <RANKING place="4" resultid="254" />
                    <RANKING place="2" resultid="593" />
                    <RANKING place="1" resultid="759" />
                    <RANKING place="3" resultid="760" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7" agemax="123" agemin="18" name="Thüringen: Kategorie I (Jg.2005 u.ä.)">
                  <RANKINGS>
                    <RANKING place="1" resultid="333" />
                    <RANKING place="2" resultid="874" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2" agemax="-1" agemin="180" easy.ak="180" calculate="TOTAL" name="Thüringen: Master I (Gesamtalter &lt;= 180 Jahre)">
                  <RANKINGS>
                    <RANKING place="1" resultid="815" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3" agemax="-1" agemin="400" easy.ak="400" calculate="TOTAL" name="Thüringen: Master II (Gesamtalter &gt; 181 Jahre)">
                  <RANKINGS>
                    <RANKING place="1" resultid="334" />
                    <RANKING place="2" resultid="816" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4" agemax="-1" agemin="400" easy.ak="400" calculate="TOTAL" name="Offene Wertung Master">
                  <RANKINGS>
                    <RANKING place="1" resultid="334" />
                    <RANKING place="3" resultid="815" />
                    <RANKING place="2" resultid="816" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8" agemax="123" agemin="1" name="Offene Wertung">
                  <RANKINGS>
                    <RANKING place="5" resultid="90" />
                    <RANKING place="2" resultid="203" />
                    <RANKING place="10" resultid="254" />
                    <RANKING place="3" resultid="333" />
                    <RANKING place="1" resultid="403" />
                    <RANKING place="9" resultid="444" />
                    <RANKING place="7" resultid="593" />
                    <RANKING place="6" resultid="759" />
                    <RANKING place="8" resultid="760" />
                    <RANKING place="4" resultid="874" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="22" number="22" gender="X" round="TIM">
              <SWIMSTYLE stroke="SURFACE" relaycount="1" distance="1500" />
              <FEE value="500" currency="EUR" />
              <HEATS>
                <HEAT heatid="22001" number="1" />
                <HEAT heatid="22002" number="2" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="9" agemin="12" name="weiblich Thüringen: Kategorie G (Jg.2014 u.j.)" />
                <AGEGROUP agegroupid="2" agemax="10" agemin="12" name="weiblich Thüringen: Kategorie F (Jg.2013)" />
                <AGEGROUP agegroupid="3" agemax="11" agemin="12" name="weiblich Thüringen: Kategorie E (Jg.2012)" />
                <AGEGROUP agegroupid="4" agemax="13" agemin="12" name="weiblich Thüringen: Kategorie D (Jg.2010/2011)" />
                <AGEGROUP agegroupid="5" agemax="15" agemin="14" name="weiblich Thüringen: Kategorie C (Jg.2008/2009)">
                  <RANKINGS>
                    <RANKING place="1" resultid="728" />
                    <RANKING place="2" resultid="905" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6" agemax="17" agemin="16" name="weiblich Thüringen: Kategorie B (Jg.2006/2007)" />
                <AGEGROUP agegroupid="7" agemax="30" agemin="18" name="weiblich Thüringen: Kategorie A (Jg.2005 u.ä.)">
                  <RANKINGS>
                    <RANKING place="1" resultid="482" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8" agemax="34" agemin="29" name="weiblich Thüringen: Master A (Jg.1989-1994)" />
                <AGEGROUP agegroupid="9" agemax="44" agemin="35" name="weiblich Thüringen: Master B (Jg.1979-1988)" />
                <AGEGROUP agegroupid="10" agemax="54" agemin="45" name="weiblich Thüringen: Master C (Jg.1969-1978)" />
                <AGEGROUP agegroupid="11" agemax="64" agemin="55" name="weiblich Thüringen: Master D (Jg.1959-1968)" />
                <AGEGROUP agegroupid="12" agemax="123" agemin="65" name="weiblich Thüringen: Master E (Jg.1958 u.ä.)" />
                <AGEGROUP agegroupid="13" agemax="123" agemin="29" name="weiblich: Offene Wertung Master" />
                <AGEGROUP agegroupid="14" agemax="30" agemin="12" name="weiblich: Offene Wertung">
                  <RANKINGS>
                    <RANKING place="2" resultid="152" />
                    <RANKING place="1" resultid="153" />
                    <RANKING place="4" resultid="198" />
                    <RANKING place="3" resultid="482" />
                    <RANKING place="5" resultid="728" />
                    <RANKING place="6" resultid="905" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="15" agemax="9" agemin="12" name="männlich Thüringen: Kategorie G (Jg.2014 u.j.)" />
                <AGEGROUP agegroupid="16" agemax="10" agemin="12" name="männlich Thüringen: Kategorie F (Jg.2013)" />
                <AGEGROUP agegroupid="17" agemax="11" agemin="12" name="männlich Thüringen: Kategorie E (Jg.2012)" />
                <AGEGROUP agegroupid="18" agemax="13" agemin="12" name="männlich Thüringen: Kategorie D (Jg.2010/2011)" />
                <AGEGROUP agegroupid="19" agemax="15" agemin="14" name="männlich Thüringen: Kategorie C (Jg.2008/2009)" />
                <AGEGROUP agegroupid="20" agemax="17" agemin="16" name="männlich Thüringen: Kategorie B (Jg.2006/2007)">
                  <RANKINGS>
                    <RANKING place="1" resultid="899" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="21" agemax="44" agemin="18" name="männlich Thüringen: Kategorie A (Jg.2005 u.ä.)" />
                <AGEGROUP agegroupid="22" agemax="34" agemin="29" name="männlich Thüringen: Master A (Jg.1989-1994)" />
                <AGEGROUP agegroupid="23" agemax="43" agemin="35" name="männlich Thüringen: Master B (Jg.1979-1988)" />
                <AGEGROUP agegroupid="24" agemax="54" agemin="45" name="männlich Thüringen: Master C (Jg.1969-1978)" />
                <AGEGROUP agegroupid="25" agemax="64" agemin="55" name="männlich Thüringen: Master D (Jg.1959-1968)" />
                <AGEGROUP agegroupid="26" agemax="123" agemin="65" name="männlich Thüringen: Master E (Jg.1958 u.ä.)" />
                <AGEGROUP agegroupid="27" agemax="123" agemin="45" name="männlich: Offene Wertung Master" />
                <AGEGROUP agegroupid="28" agemax="44" agemin="12" name="männlich: Offene Wertung">
                  <RANKINGS>
                    <RANKING place="1" resultid="47" />
                    <RANKING place="2" resultid="899" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
          </EVENTS>
        </SESSION>
      </SESSIONS>
      <CLUBS>
        <CLUB name="1. Chemnitzer Tauchverein e.V." nation="GER" region="20" code="0">
          <ATHLETES>
            <ATHLETE athleteid="168" birthdate="2005-01-01" gender="M" lastname="Porges" firstname="Marcel" license="0">
              <RESULTS>
                <RESULT resultid="527" eventid="2" swimtime="00:00:16.52" lane="4" heatid="2005" />
                <RESULT resultid="528" eventid="7" swimtime="00:07:13.98" lane="4" heatid="7004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:49.45" />
                    <SPLIT distance="200" swimtime="00:01:42.70" />
                    <SPLIT distance="300" swimtime="00:02:38.20" />
                    <SPLIT distance="400" swimtime="00:03:34.44" />
                    <SPLIT distance="500" swimtime="00:04:30.63" />
                    <SPLIT distance="600" swimtime="00:05:26.43" />
                    <SPLIT distance="700" swimtime="00:06:21.98" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="529" eventid="17" swimtime="00:03:26.93" lane="5" heatid="17004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:47.61" />
                    <SPLIT distance="200" swimtime="00:01:41.29" />
                    <SPLIT distance="300" swimtime="00:02:34.76" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="530" eventid="19" swimtime="00:00:39.50" lane="6" heatid="19004" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="169" birthdate="2006-01-01" gender="M" lastname="Lorenz" firstname="Emil" license="0">
              <RESULTS>
                <RESULT resultid="531" eventid="2" swimtime="00:00:17.63" lane="2" heatid="2006" />
                <RESULT resultid="532" eventid="9" status="DSQ" swimtime="00:00:00.00" lane="5" heatid="9009" comment="aufgegeben nach 18m" />
                <RESULT resultid="533" eventid="12" swimtime="00:00:19.97" lane="5" heatid="12008" />
                <RESULT resultid="534" eventid="19" swimtime="00:00:44.14" lane="8" heatid="19004" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="170" birthdate="2007-01-01" gender="F" lastname="Ullrich" firstname="Johanna Hermine" license="0">
              <RESULTS>
                <RESULT resultid="535" eventid="1" swimtime="00:00:24.77" lane="8" heatid="1004" />
                <RESULT resultid="536" eventid="8" swimtime="00:00:56.34" lane="3" heatid="8011" />
                <RESULT resultid="537" eventid="11" swimtime="00:00:25.79" lane="3" heatid="11011" />
                <RESULT resultid="538" eventid="18" swimtime="00:00:58.29" lane="6" heatid="18003" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="171" birthdate="2008-01-01" gender="F" lastname="Franke" firstname="Jenny" license="0">
              <RESULTS>
                <RESULT resultid="539" eventid="1" swimtime="00:00:22.47" lane="7" heatid="1005" />
                <RESULT resultid="540" eventid="8" swimtime="00:00:54.10" lane="8" heatid="8012" />
                <RESULT resultid="541" eventid="11" swimtime="00:00:24.59" lane="6" heatid="11012" />
                <RESULT resultid="542" eventid="16" swimtime="00:04:49.05" lane="4" heatid="16005">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:03.13" />
                    <SPLIT distance="200" swimtime="00:02:15.47" />
                    <SPLIT distance="300" swimtime="00:03:33.12" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="172" birthdate="2009-01-01" gender="M" lastname="Hans" firstname="Yannick" license="0">
              <RESULTS>
                <RESULT resultid="543" eventid="2" swimtime="00:00:24.44" lane="2" heatid="2002" />
                <RESULT resultid="544" eventid="9" swimtime="00:00:55.36" lane="3" heatid="9006" />
                <RESULT resultid="545" eventid="12" swimtime="00:00:24.75" lane="2" heatid="12006" />
                <RESULT resultid="546" eventid="17" swimtime="00:04:21.45" lane="4" heatid="17002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:58.11" />
                    <SPLIT distance="200" swimtime="00:02:08.24" />
                    <SPLIT distance="300" swimtime="00:03:18.91" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="173" birthdate="2010-01-01" gender="F" lastname="Schwarzer" firstname="Angelina Sophie" license="0">
              <RESULTS>
                <RESULT resultid="547" eventid="3" swimtime="00:00:29.85" lane="6" heatid="3001" />
                <RESULT resultid="548" eventid="8" swimtime="00:00:58.40" lane="8" heatid="8010" />
                <RESULT resultid="549" eventid="11" swimtime="00:00:26.20" lane="5" heatid="11008" />
                <RESULT resultid="550" eventid="16" swimtime="00:04:56.13" lane="2" heatid="16005">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:07.67" />
                    <SPLIT distance="200" swimtime="00:02:25.45" />
                    <SPLIT distance="300" swimtime="00:03:45.44" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="174" birthdate="2011-01-01" gender="F" lastname="Nisch" firstname="Hanna Maria" license="0">
              <RESULTS>
                <RESULT resultid="551" eventid="3" status="DSQ" swimtime="00:00:44.21" lane="3" heatid="3001" comment="Gesicht aus dem Wasser bei 20m" />
                <RESULT resultid="552" eventid="8" swimtime="00:01:01.18" lane="4" heatid="8008" />
                <RESULT resultid="553" eventid="11" swimtime="00:00:27.00" lane="6" heatid="11008" />
                <RESULT resultid="554" eventid="16" swimtime="00:04:55.03" lane="5" heatid="16004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:10.49" />
                    <SPLIT distance="200" swimtime="00:02:28.17" />
                    <SPLIT distance="300" swimtime="00:03:45.82" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="Aquanauten Karlsruhe-Durlach e.V." nation="GER" region="33" code="0">
          <ATHLETES>
            <ATHLETE athleteid="29" birthdate="2007-01-01" gender="F" lastname="Haag" firstname="Jenny" license="0">
              <RESULTS>
                <RESULT resultid="117" eventid="1" swimtime="00:00:28.99" lane="3" heatid="1001" />
                <RESULT resultid="113" eventid="8" swimtime="00:01:06.87" lane="3" heatid="8004" />
                <RESULT resultid="119" eventid="11" swimtime="00:00:30.25" lane="2" heatid="11006" />
                <RESULT resultid="115" eventid="13" swimtime="00:02:37.12" lane="3" heatid="13003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:12.37" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="30" birthdate="2007-01-01" gender="F" lastname="Kirchner" firstname="Nia" license="0">
              <RESULTS>
                <RESULT resultid="116" eventid="1" swimtime="00:00:24.31" lane="6" heatid="1003" />
                <RESULT resultid="120" eventid="7" status="DSQ" swimtime="00:00:00.00" lane="1" heatid="7002" comment="aufgegeben nach 140m">
                  <SPLITS>
                    <SPLIT distance="200" swimtime="00:01:04.08" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="118" eventid="11" swimtime="00:00:24.76" lane="7" heatid="11009" />
                <RESULT resultid="114" eventid="18" swimtime="00:00:57.11" lane="3" heatid="18002" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="Berliner TSC e.V." nation="GER" region="21" code="0">
          <ATHLETES>
            <ATHLETE athleteid="1" birthdate="2007-01-01" gender="F" lastname="Manthey" firstname="Maxime" license="0">
              <RESULTS>
                <RESULT resultid="24" eventid="1" swimtime="00:00:17.71" lane="2" heatid="1007" />
                <RESULT resultid="1" eventid="8" swimtime="00:00:47.10" lane="2" heatid="8014" />
                <RESULT resultid="32" eventid="11" swimtime="00:00:20.35" lane="6" heatid="11014" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="2" birthdate="2007-01-01" gender="F" lastname="Eggert" firstname="Emilia" license="0">
              <RESULTS>
                <RESULT resultid="25" eventid="1" swimtime="00:00:18.85" lane="6" heatid="1006" />
                <RESULT resultid="2" eventid="8" swimtime="00:00:45.05" lane="1" heatid="8014" />
                <RESULT resultid="10" eventid="13" swimtime="00:01:44.00" lane="6" heatid="13011">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:50.85" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="17" eventid="16" swimtime="00:03:47.82" lane="4" heatid="16007">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:52.03" />
                    <SPLIT distance="200" swimtime="00:01:51.10" />
                    <SPLIT distance="300" swimtime="00:02:51.16" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="3" birthdate="2008-01-01" gender="F" lastname="Bublitz" firstname="Tessa" license="0">
              <RESULTS>
                <RESULT resultid="27" eventid="1" swimtime="00:00:19.79" lane="6" heatid="1004" />
                <RESULT resultid="3" eventid="8" swimtime="00:00:47.78" lane="3" heatid="8012" />
                <RESULT resultid="11" eventid="13" swimtime="00:01:47.59" lane="1" heatid="13010">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:52.26" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="18" eventid="16" swimtime="00:03:52.35" lane="6" heatid="16006">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:53.30" />
                    <SPLIT distance="200" swimtime="00:01:53.54" />
                    <SPLIT distance="300" swimtime="00:02:54.83" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="4" birthdate="2007-01-01" gender="F" lastname="Beske" firstname="Lena" license="0">
              <RESULTS>
                <RESULT resultid="26" eventid="1" swimtime="00:00:21.70" lane="5" heatid="1004" />
                <RESULT resultid="4" eventid="8" swimtime="00:00:56.84" lane="5" heatid="8010" />
                <RESULT resultid="33" eventid="11" swimtime="00:00:23.00" lane="1" heatid="11012" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="5" birthdate="2005-01-01" gender="F" lastname="Seidler" firstname="Anika" license="0">
              <RESULTS>
                <RESULT resultid="28" eventid="1" swimtime="00:00:25.00" lane="4" heatid="1003" />
                <RESULT resultid="5" eventid="8" swimtime="00:01:00.32" lane="2" heatid="8009" />
                <RESULT resultid="35" eventid="11" swimtime="00:00:27.44" lane="4" heatid="11008" />
                <RESULT resultid="12" eventid="13" swimtime="00:02:13.50" lane="8" heatid="13008">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:02.94" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="6" birthdate="2011-01-01" gender="F" lastname="Stobbe" firstname="Bella" license="0">
              <RESULTS>
                <RESULT resultid="6" eventid="8" swimtime="00:01:00.90" lane="8" heatid="8009" />
                <RESULT resultid="34" eventid="11" swimtime="00:00:26.65" lane="7" heatid="11011" />
                <RESULT resultid="13" eventid="13" swimtime="00:02:12.46" lane="6" heatid="13006">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:03.72" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="19" eventid="16" status="DNS" swimtime="00:00:00.00" lane="3" heatid="16003" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="7" birthdate="2008-01-01" gender="M" lastname="Welke" firstname="Anton" license="0">
              <RESULTS>
                <RESULT resultid="30" eventid="2" swimtime="00:00:18.70" lane="1" heatid="2005" />
                <RESULT resultid="7" eventid="9" swimtime="00:00:46.02" lane="2" heatid="9009" />
                <RESULT resultid="15" eventid="14" swimtime="00:01:41.32" lane="6" heatid="14006">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:49.63" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="20" eventid="17" swimtime="00:03:45.00" lane="2" heatid="17004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:50.88" />
                    <SPLIT distance="200" swimtime="00:01:49.22" />
                    <SPLIT distance="300" swimtime="00:02:48.03" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="8" birthdate="2009-01-01" gender="M" lastname="Martiny" firstname="Peter" license="0">
              <RESULTS>
                <RESULT resultid="31" eventid="2" swimtime="00:00:20.97" lane="5" heatid="2002" />
                <RESULT resultid="8" eventid="9" swimtime="00:00:51.36" lane="1" heatid="9007" />
                <RESULT resultid="16" eventid="14" swimtime="00:01:56.20" lane="1" heatid="14005">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:55.61" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="21" eventid="17" swimtime="00:04:10.00" lane="5" heatid="17003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:57.10" />
                    <SPLIT distance="200" swimtime="00:02:02.25" />
                    <SPLIT distance="300" swimtime="00:03:08.50" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="9" birthdate="2004-01-01" gender="M" lastname="Beske" firstname="Tom" license="0">
              <RESULTS>
                <RESULT resultid="29" eventid="2" swimtime="00:00:17.28" lane="8" heatid="2006" />
                <RESULT resultid="22" eventid="10" swimtime="00:03:07.96" lane="5" heatid="10003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:44.88" />
                    <SPLIT distance="200" swimtime="00:01:33.08" />
                    <SPLIT distance="300" swimtime="00:02:22.49" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="14" eventid="14" swimtime="00:01:34.77" lane="3" heatid="14006">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:43.71" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="9" eventid="19" swimtime="00:00:38.42" lane="5" heatid="19004" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY number="1" gender="F" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="23" eventid="20" swimtime="00:03:12.19" lane="3" heatid="20003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:47.15" />
                    <SPLIT distance="200" swimtime="00:01:33.74" />
                    <SPLIT distance="300" swimtime="00:02:27.46" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1" number="1" />
                    <RELAYPOSITION athleteid="3" number="2" />
                    <RELAYPOSITION athleteid="4" number="3" />
                    <RELAYPOSITION athleteid="2" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB name="Binger Tauchsportclub e.V." nation="GER" region="29" code="0">
          <ATHLETES>
            <ATHLETE athleteid="11" birthdate="2008-01-01" gender="M" lastname="Funke" firstname="Paul" license="0">
              <RESULTS>
                <RESULT resultid="41" eventid="2" swimtime="00:00:24.42" lane="1" heatid="2002" />
                <RESULT resultid="36" eventid="9" swimtime="00:00:55.95" lane="6" heatid="9006" />
                <RESULT resultid="43" eventid="12" swimtime="00:00:25.14" lane="4" heatid="12005" />
                <RESULT resultid="39" eventid="17" swimtime="00:04:26.58" lane="3" heatid="17003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:59.83" />
                    <SPLIT distance="200" swimtime="00:02:09.63" />
                    <SPLIT distance="300" swimtime="00:03:19.27" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="47" eventid="22" swimtime="00:18:01.15" lane="2" heatid="22002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:02.17" />
                    <SPLIT distance="200" swimtime="00:02:12.06" />
                    <SPLIT distance="300" swimtime="00:03:24.12" />
                    <SPLIT distance="400" swimtime="00:04:36.35" />
                    <SPLIT distance="500" swimtime="00:05:48.58" />
                    <SPLIT distance="600" swimtime="00:06:59.29" />
                    <SPLIT distance="700" swimtime="00:08:11.12" />
                    <SPLIT distance="800" swimtime="00:09:23.17" />
                    <SPLIT distance="900" swimtime="00:10:36.40" />
                    <SPLIT distance="1000" swimtime="00:11:51.30" />
                    <SPLIT distance="1100" swimtime="00:13:07.19" />
                    <SPLIT distance="1200" swimtime="00:14:20.97" />
                    <SPLIT distance="1300" swimtime="00:15:34.55" />
                    <SPLIT distance="1400" swimtime="00:16:47.46" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="12" birthdate="2009-01-01" gender="M" lastname="Moritz" firstname="Silas" license="0">
              <RESULTS>
                <RESULT resultid="42" eventid="2" swimtime="00:00:22.84" lane="3" heatid="2001" />
                <RESULT resultid="46" eventid="7" swimtime="00:09:54.00" lane="4" heatid="7001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:05.20" />
                    <SPLIT distance="200" swimtime="00:02:17.91" />
                    <SPLIT distance="300" swimtime="00:03:32.32" />
                    <SPLIT distance="400" swimtime="00:04:50.52" />
                    <SPLIT distance="500" swimtime="00:06:09.08" />
                    <SPLIT distance="600" swimtime="00:07:26.21" />
                    <SPLIT distance="700" swimtime="00:08:39.46" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="37" eventid="9" swimtime="00:00:57.03" lane="1" heatid="9006" />
                <RESULT resultid="44" eventid="12" swimtime="00:00:27.37" lane="2" heatid="12004" />
                <RESULT resultid="38" eventid="14" swimtime="00:02:10.75" lane="6" heatid="14004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:04.17" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="40" eventid="17" swimtime="00:04:47.44" lane="5" heatid="17002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:06.81" />
                    <SPLIT distance="200" swimtime="00:02:20.24" />
                    <SPLIT distance="300" swimtime="00:03:35.01" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="KP Pardubice" nation="CZE" region="0" code="0">
          <ATHLETES>
            <ATHLETE athleteid="55" birthdate="2006-01-01" gender="F" lastname="Stránská" firstname="Tereza" license="0">
              <RESULTS>
                <RESULT resultid="192" eventid="8" swimtime="00:00:56.46" lane="2" heatid="8010" />
                <RESULT resultid="208" eventid="11" swimtime="00:00:24.72" lane="4" heatid="11010" />
                <RESULT resultid="200" eventid="16" swimtime="00:04:38.85" lane="2" heatid="16004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:06.54" />
                    <SPLIT distance="200" swimtime="00:02:17.96" />
                    <SPLIT distance="300" swimtime="00:03:30.35" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="56" birthdate="2007-01-01" gender="M" lastname="Pošva" firstname="Lukáš" license="0">
              <RESULTS>
                <RESULT resultid="207" eventid="2" swimtime="00:00:20.96" lane="3" heatid="2003" />
                <RESULT resultid="193" eventid="9" swimtime="00:00:48.48" lane="1" heatid="9008" />
                <RESULT resultid="210" eventid="12" swimtime="00:00:21.44" lane="7" heatid="12007" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="57" birthdate="2007-01-01" gender="M" lastname="Malý" firstname="Václav" license="0">
              <RESULTS>
                <RESULT resultid="206" eventid="2" swimtime="00:00:18.37" lane="4" heatid="2003" />
                <RESULT resultid="194" eventid="9" swimtime="00:00:50.53" lane="7" heatid="9007" />
                <RESULT resultid="211" eventid="12" status="DSQ" swimtime="00:00:21.23" lane="5" heatid="12006" comment="15m nach Start übertaucht" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="58" birthdate="2006-01-01" gender="F" lastname="Koryntová" firstname="Alžbìta" license="0">
              <RESULTS>
                <RESULT resultid="215" eventid="7" swimtime="00:08:30.47" lane="3" heatid="7003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:56.16" />
                    <SPLIT distance="200" swimtime="00:01:57.13" />
                    <SPLIT distance="300" swimtime="00:02:59.31" />
                    <SPLIT distance="400" swimtime="00:04:04.38" />
                    <SPLIT distance="500" swimtime="00:05:10.86" />
                    <SPLIT distance="600" swimtime="00:06:18.34" />
                    <SPLIT distance="700" swimtime="00:07:25.49" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="214" eventid="13" swimtime="00:01:53.78" lane="4" heatid="13009">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:53.51" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="195" eventid="18" swimtime="00:00:47.92" lane="7" heatid="18004" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="59" birthdate="2007-01-01" gender="F" lastname="Malá" firstname="Lea" license="0">
              <RESULTS>
                <RESULT resultid="202" eventid="10" swimtime="00:04:13.16" lane="2" heatid="10002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:57.34" />
                    <SPLIT distance="200" swimtime="00:02:02.82" />
                    <SPLIT distance="300" swimtime="00:03:10.59" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="196" eventid="18" swimtime="00:00:49.16" lane="4" heatid="18003" />
                <RESULT resultid="198" eventid="22" swimtime="00:18:15.71" lane="6" heatid="22001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:05.53" />
                    <SPLIT distance="200" swimtime="00:02:15.81" />
                    <SPLIT distance="300" swimtime="00:03:28.69" />
                    <SPLIT distance="400" swimtime="00:04:41.67" />
                    <SPLIT distance="500" swimtime="00:05:54.29" />
                    <SPLIT distance="600" swimtime="00:07:06.96" />
                    <SPLIT distance="700" swimtime="00:08:21.08" />
                    <SPLIT distance="800" swimtime="00:09:36.57" />
                    <SPLIT distance="900" swimtime="00:10:50.58" />
                    <SPLIT distance="1000" swimtime="00:12:05.24" />
                    <SPLIT distance="1100" swimtime="00:13:21.16" />
                    <SPLIT distance="1200" swimtime="00:14:37.41" />
                    <SPLIT distance="1300" swimtime="00:15:54.37" />
                    <SPLIT distance="1400" swimtime="00:17:08.26" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="60" birthdate="2004-01-01" gender="M" lastname="Cimburek" firstname="Daniel" license="0">
              <RESULTS>
                <RESULT resultid="204" eventid="2" swimtime="00:00:17.09" lane="6" heatid="2006" />
                <RESULT resultid="201" eventid="10" swimtime="00:03:07.31" lane="4" heatid="10003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:45.06" />
                    <SPLIT distance="200" swimtime="00:01:33.36" />
                    <SPLIT distance="300" swimtime="00:02:21.13" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="197" eventid="19" swimtime="00:00:36.29" lane="4" heatid="19004" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="63" birthdate="2003-01-01" gender="M" lastname="Kvìton" firstname="Jan" license="0">
              <RESULTS>
                <RESULT resultid="205" eventid="2" status="DSQ" swimtime="00:00:00.00" lane="7" heatid="2006" comment="Gesicht aus dem Wasser bei 40m" />
                <RESULT resultid="213" eventid="12" swimtime="00:00:19.82" lane="4" heatid="12008" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY number="1" gender="M" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="203" eventid="21" swimtime="00:03:00.41" lane="3" heatid="21002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:44.72" />
                    <SPLIT distance="200" swimtime="00:01:31.93" />
                    <SPLIT distance="300" swimtime="00:02:20.71" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="63" number="1" />
                    <RELAYPOSITION athleteid="56" number="2" />
                    <RELAYPOSITION athleteid="57" number="3" />
                    <RELAYPOSITION athleteid="60" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB name="SC DHfK Leipzig Flossenschwimmen" nation="GER" region="20" code="0">
          <ATHLETES>
            <ATHLETE athleteid="120" birthdate="2008-01-01" gender="F" lastname="Horenok" firstname="Maiia" license="0">
              <RESULTS>
                <RESULT resultid="404" eventid="1" swimtime="00:00:18.51" lane="1" heatid="1006" />
                <RESULT resultid="379" eventid="8" swimtime="00:00:45.55" lane="6" heatid="8013" />
                <RESULT resultid="407" eventid="11" swimtime="00:00:20.01" lane="2" heatid="11014" />
                <RESULT resultid="394" eventid="16" swimtime="00:03:48.49" lane="7" heatid="16007">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:53.68" />
                    <SPLIT distance="200" swimtime="00:01:53.26" />
                    <SPLIT distance="300" swimtime="00:02:53.31" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="121" birthdate="2008-01-01" gender="F" lastname="Kulchytska" firstname="Polina" license="0">
              <RESULTS>
                <RESULT resultid="380" eventid="8" swimtime="00:00:49.61" lane="5" heatid="8012" />
                <RESULT resultid="391" eventid="13" swimtime="00:01:50.68" lane="5" heatid="13009">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:53.81" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="395" eventid="16" swimtime="00:03:54.78" lane="1" heatid="16007">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:54.94" />
                    <SPLIT distance="200" swimtime="00:01:55.18" />
                    <SPLIT distance="300" swimtime="00:02:56.07" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="387" eventid="18" swimtime="00:00:47.45" lane="6" heatid="18004" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="123" birthdate="2001-01-01" gender="M" lastname="Mörstedt" firstname="Justus" license="0">
              <RESULTS>
                <RESULT resultid="382" eventid="9" swimtime="00:00:35.42" lane="4" heatid="9010" />
                <RESULT resultid="392" eventid="14" swimtime="00:01:22.46" lane="4" heatid="14006">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:40.01" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="124" birthdate="2001-01-01" gender="M" lastname="Gaida" firstname="Duncan" license="0">
              <RESULTS>
                <RESULT resultid="383" eventid="9" swimtime="00:00:37.54" lane="3" heatid="9010" />
                <RESULT resultid="398" eventid="17" swimtime="00:03:15.19" lane="4" heatid="17004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:46.10" />
                    <SPLIT distance="200" swimtime="00:01:35.65" />
                    <SPLIT distance="300" swimtime="00:02:25.89" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="125" birthdate="1999-01-01" gender="M" lastname="Wahlstadt" firstname="Felix" license="0">
              <RESULTS>
                <RESULT resultid="384" eventid="9" swimtime="00:00:40.01" lane="2" heatid="9010" />
                <RESULT resultid="409" eventid="12" swimtime="00:00:17.98" lane="3" heatid="12009" />
                <RESULT resultid="399" eventid="17" swimtime="00:03:27.71" lane="6" heatid="17004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:48.34" />
                    <SPLIT distance="200" swimtime="00:01:42.15" />
                    <SPLIT distance="300" swimtime="00:02:36.09" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="126" birthdate="2009-01-01" gender="M" lastname="Batiuk" firstname="Mykyta" license="0">
              <RESULTS>
                <RESULT resultid="405" eventid="2" swimtime="00:00:19.04" lane="5" heatid="2005" />
                <RESULT resultid="385" eventid="9" swimtime="00:00:47.77" lane="1" heatid="9010" />
                <RESULT resultid="410" eventid="12" swimtime="00:00:20.40" lane="2" heatid="12009" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="127" birthdate="2008-01-01" gender="M" lastname="Berger" firstname="Alex Michael" license="0">
              <RESULTS>
                <RESULT resultid="386" eventid="9" swimtime="00:00:50.32" lane="3" heatid="9007" />
                <RESULT resultid="412" eventid="12" swimtime="00:00:22.83" lane="1" heatid="12007" />
                <RESULT resultid="401" eventid="17" swimtime="00:04:07.62" lane="4" heatid="17003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:56.51" />
                    <SPLIT distance="200" swimtime="00:02:02.03" />
                    <SPLIT distance="300" swimtime="00:03:07.86" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="128" birthdate="2007-01-01" gender="F" lastname="Holtz" firstname="Leonie-Florentine" license="0">
              <RESULTS>
                <RESULT resultid="408" eventid="11" swimtime="00:00:22.77" lane="4" heatid="11012" />
                <RESULT resultid="396" eventid="16" swimtime="00:04:13.23" lane="3" heatid="16006">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:58.23" />
                    <SPLIT distance="200" swimtime="00:02:03.73" />
                    <SPLIT distance="300" swimtime="00:03:09.74" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="388" eventid="18" swimtime="00:00:50.75" lane="8" heatid="18004" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="129" birthdate="2007-01-01" gender="F" lastname="Hempler" firstname="Emily" license="0">
              <RESULTS>
                <RESULT resultid="413" eventid="7" swimtime="00:07:37.78" lane="5" heatid="7004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:51.68" />
                    <SPLIT distance="200" swimtime="00:01:48.92" />
                    <SPLIT distance="300" swimtime="00:02:46.45" />
                    <SPLIT distance="400" swimtime="00:03:44.98" />
                    <SPLIT distance="500" swimtime="00:04:43.30" />
                    <SPLIT distance="600" swimtime="00:05:42.00" />
                    <SPLIT distance="700" swimtime="00:06:40.74" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="390" eventid="13" swimtime="00:01:43.15" lane="2" heatid="13011">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:49.49" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="393" eventid="16" swimtime="00:03:38.72" lane="5" heatid="16008">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:51.16" />
                    <SPLIT distance="200" swimtime="00:01:46.36" />
                    <SPLIT distance="300" swimtime="00:02:42.58" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="307" birthdate="1984-01-01" gender="F" lastname="Sapsai" firstname="Irina" license="0">
              <RESULTS>
                <RESULT resultid="956" eventid="11" swimtime="00:00:25.76" lane="2" heatid="11011" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="308" birthdate="1977-01-01" gender="M" lastname="Nehrdich" firstname="Thomas" license="0">
              <RESULTS>
                <RESULT resultid="957" eventid="9" swimtime="00:00:47.48" lane="3" heatid="9008" />
                <RESULT resultid="958" eventid="12" swimtime="00:00:20.52" lane="3" heatid="12007" />
                <RESULT resultid="959" eventid="14" swimtime="00:01:49.26" lane="5" heatid="14005">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:52.29" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="960" eventid="17" swimtime="00:04:02.68" lane="7" heatid="17004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:54.22" />
                    <SPLIT distance="200" swimtime="00:01:55.99" />
                    <SPLIT distance="300" swimtime="00:03:01.73" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY number="1" gender="F" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="402" eventid="20" swimtime="00:03:11.51" lane="4" heatid="20003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:46.74" />
                    <SPLIT distance="200" swimtime="00:01:36.23" />
                    <SPLIT distance="300" swimtime="00:02:27.32" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="129" number="1" />
                    <RELAYPOSITION athleteid="121" number="2" />
                    <RELAYPOSITION athleteid="128" number="3" />
                    <RELAYPOSITION athleteid="120" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" gender="M" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="403" eventid="21" swimtime="00:02:57.25" lane="5" heatid="21002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:40.81" />
                    <SPLIT distance="200" swimtime="00:01:28.20" />
                    <SPLIT distance="300" swimtime="00:02:18.65" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="125" number="1" />
                    <RELAYPOSITION athleteid="126" number="2" />
                    <RELAYPOSITION athleteid="127" number="3" />
                    <RELAYPOSITION athleteid="124" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB name="SC Riesa Sekt. Flossenschwimmen" nation="GER" region="20" code="0">
          <ATHLETES>
            <ATHLETE athleteid="13" birthdate="2006-01-01" gender="M" lastname="Loßner" firstname="Niklas" license="0">
              <RESULTS>
                <RESULT resultid="50" eventid="2" swimtime="00:00:15.34" lane="4" heatid="2006" />
                <RESULT resultid="48" eventid="9" swimtime="00:00:38.76" lane="6" heatid="9010" />
                <RESULT resultid="51" eventid="12" swimtime="00:00:16.71" lane="5" heatid="12009" />
                <RESULT resultid="49" eventid="17" swimtime="00:03:32.82" lane="3" heatid="17004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:46.42" />
                    <SPLIT distance="200" swimtime="00:01:41.17" />
                    <SPLIT distance="300" swimtime="00:02:38.60" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="SG Dresden" nation="GER" region="20" code="0">
          <ATHLETES>
            <ATHLETE athleteid="216" birthdate="1986-01-01" gender="F" lastname="Klar" firstname="Margarethe" license="0">
              <RESULTS>
                <RESULT resultid="675" eventid="1" swimtime="00:00:26.46" lane="7" heatid="1003" />
                <RESULT resultid="676" eventid="8" swimtime="00:01:00.41" lane="6" heatid="8010" />
                <RESULT resultid="677" eventid="11" swimtime="00:00:28.26" lane="8" heatid="11010" />
                <RESULT resultid="678" eventid="18" swimtime="00:00:58.97" lane="3" heatid="18003" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="217" birthdate="2000-01-01" gender="F" lastname="Rütze" firstname="Michel" license="0">
              <RESULTS>
                <RESULT resultid="679" eventid="1" swimtime="00:00:17.14" lane="4" heatid="1007" />
                <RESULT resultid="680" eventid="8" swimtime="00:00:41.16" lane="4" heatid="8014" />
                <RESULT resultid="681" eventid="13" swimtime="00:01:33.63" lane="4" heatid="13011">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:44.80" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="682" eventid="18" swimtime="00:00:39.80" lane="4" heatid="18005" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="218" birthdate="2004-01-01" gender="F" lastname="Placzek" firstname="Lilly" license="0">
              <RESULTS>
                <RESULT resultid="683" eventid="1" swimtime="00:00:17.79" lane="3" heatid="1007" />
                <RESULT resultid="684" eventid="8" swimtime="00:00:44.88" lane="7" heatid="8014" />
                <RESULT resultid="685" eventid="13" swimtime="00:01:44.13" lane="8" heatid="13011">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:48.99" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="686" eventid="18" swimtime="00:00:41.72" lane="3" heatid="18005" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="219" birthdate="2005-01-01" gender="F" lastname="Richter" firstname="Franca" license="0">
              <RESULTS>
                <RESULT resultid="687" eventid="10" status="DNS" swimtime="00:00:00.00" lane="6" heatid="10003" />
                <RESULT resultid="688" eventid="13" swimtime="00:02:02.67" lane="7" heatid="13011">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:58.25" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="689" eventid="16" swimtime="00:04:27.38" lane="2" heatid="16008">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:03.06" />
                    <SPLIT distance="200" swimtime="00:02:11.86" />
                    <SPLIT distance="300" swimtime="00:03:20.25" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="690" eventid="18" status="DNS" swimtime="00:00:00.00" lane="2" heatid="18005" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="SG Finswimming Jena" nation="GER" region="35" code="0">
          <ATHLETES>
            <ATHLETE athleteid="151" birthdate="1979-01-01" gender="M" lastname="Schubert" firstname="Michael" license="0">
              <RESULTS>
                <RESULT resultid="471" eventid="10" swimtime="00:06:25.49" lane="3" heatid="10001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:22.13" />
                    <SPLIT distance="200" swimtime="00:03:02.13" />
                    <SPLIT distance="300" swimtime="00:04:42.97" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="472" eventid="19" swimtime="00:01:13.79" lane="4" heatid="19001" />
                <RESULT resultid="473" eventid="22" status="DSQ" swimtime="00:00:00.00" lane="7" heatid="22001" comment="aufgegeben nach 300m" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="152" birthdate="1999-01-01" gender="F" lastname="Jacke" firstname="Lena" license="0">
              <RESULTS>
                <RESULT resultid="474" eventid="7" swimtime="00:08:52.16" lane="8" heatid="7003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:02.86" />
                    <SPLIT distance="200" swimtime="00:02:07.77" />
                    <SPLIT distance="300" swimtime="00:03:16.19" />
                    <SPLIT distance="400" swimtime="00:04:23.36" />
                    <SPLIT distance="500" swimtime="00:05:33.83" />
                    <SPLIT distance="600" swimtime="00:06:41.55" />
                    <SPLIT distance="700" swimtime="00:07:51.17" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="475" eventid="10" swimtime="00:04:26.43" lane="1" heatid="10002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:01.09" />
                    <SPLIT distance="200" swimtime="00:02:08.02" />
                    <SPLIT distance="300" swimtime="00:03:20.00" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="476" eventid="16" swimtime="00:04:12.27" lane="2" heatid="16006">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:01.75" />
                    <SPLIT distance="200" swimtime="00:02:05.67" />
                    <SPLIT distance="300" swimtime="00:03:10.78" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="154" birthdate="2005-01-01" gender="F" lastname="Altenstein" firstname="Louise" license="0">
              <RESULTS>
                <RESULT resultid="478" eventid="7" swimtime="00:08:26.28" lane="1" heatid="7004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:58.16" />
                    <SPLIT distance="200" swimtime="00:02:00.07" />
                    <SPLIT distance="300" swimtime="00:03:03.98" />
                    <SPLIT distance="400" swimtime="00:04:08.02" />
                    <SPLIT distance="500" swimtime="00:05:12.73" />
                    <SPLIT distance="600" swimtime="00:06:18.15" />
                    <SPLIT distance="700" swimtime="00:07:24.20" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="479" eventid="10" swimtime="00:04:01.23" lane="6" heatid="10002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:55.00" />
                    <SPLIT distance="200" swimtime="00:01:57.56" />
                    <SPLIT distance="300" swimtime="00:03:01.05" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="480" eventid="16" swimtime="00:03:57.31" lane="6" heatid="16007">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:55.41" />
                    <SPLIT distance="200" swimtime="00:01:56.38" />
                    <SPLIT distance="300" swimtime="00:02:58.42" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="481" eventid="18" swimtime="00:00:46.67" lane="3" heatid="18004" />
                <RESULT resultid="482" eventid="22" swimtime="00:17:18.00" lane="6" heatid="22002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:04.81" />
                    <SPLIT distance="200" swimtime="00:02:12.83" />
                    <SPLIT distance="300" swimtime="00:03:22.32" />
                    <SPLIT distance="400" swimtime="00:04:31.53" />
                    <SPLIT distance="500" swimtime="00:05:40.96" />
                    <SPLIT distance="600" swimtime="00:06:50.83" />
                    <SPLIT distance="700" swimtime="00:08:01.32" />
                    <SPLIT distance="800" swimtime="00:09:11.66" />
                    <SPLIT distance="900" swimtime="00:10:20.98" />
                    <SPLIT distance="1000" swimtime="00:11:31.08" />
                    <SPLIT distance="1100" swimtime="00:12:40.63" />
                    <SPLIT distance="1200" swimtime="00:13:49.09" />
                    <SPLIT distance="1300" swimtime="00:15:00.27" />
                    <SPLIT distance="1400" swimtime="00:16:10.65" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="155" birthdate="2005-01-01" gender="M" lastname="Preuß" firstname="Marek" license="0">
              <RESULTS>
                <RESULT resultid="483" eventid="7" status="DNS" swimtime="00:00:00.00" lane="4" heatid="7003" />
                <RESULT resultid="484" eventid="10" status="DNS" swimtime="00:00:00.00" lane="5" heatid="10002" />
                <RESULT resultid="485" eventid="17" status="DNS" swimtime="00:00:00.00" lane="1" heatid="17004" />
                <RESULT resultid="486" eventid="19" status="DNS" swimtime="00:00:00.00" lane="1" heatid="19003" />
                <RESULT resultid="487" eventid="22" status="DNS" swimtime="00:00:00.00" lane="3" heatid="22002" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="157" birthdate="2006-01-01" gender="F" lastname="Fabian" firstname="Lareen" license="0">
              <RESULTS>
                <RESULT resultid="489" eventid="1" swimtime="00:00:22.88" lane="2" heatid="1004" />
                <RESULT resultid="490" eventid="7" swimtime="00:10:15.56" lane="2" heatid="7002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:04.37" />
                    <SPLIT distance="200" swimtime="00:02:18.07" />
                    <SPLIT distance="300" swimtime="00:03:34.68" />
                    <SPLIT distance="400" swimtime="00:04:55.30" />
                    <SPLIT distance="500" swimtime="00:06:16.52" />
                    <SPLIT distance="600" swimtime="00:07:40.38" />
                    <SPLIT distance="700" swimtime="00:09:00.57" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="491" eventid="11" swimtime="00:00:25.70" lane="6" heatid="11011" />
                <RESULT resultid="492" eventid="13" swimtime="00:02:09.65" lane="1" heatid="13008">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:01.83" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="493" eventid="18" swimtime="00:01:02.15" lane="7" heatid="18003" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="158" birthdate="2006-01-01" gender="F" lastname="Steininger" firstname="Liese" license="0">
              <RESULTS>
                <RESULT resultid="494" eventid="7" swimtime="00:10:46.25" lane="5" heatid="7001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:13.50" />
                    <SPLIT distance="200" swimtime="00:02:34.84" />
                    <SPLIT distance="300" swimtime="00:03:52.80" />
                    <SPLIT distance="400" swimtime="00:05:20.61" />
                    <SPLIT distance="500" swimtime="00:06:47.32" />
                    <SPLIT distance="600" swimtime="00:08:06.75" />
                    <SPLIT distance="700" swimtime="00:09:31.83" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="495" eventid="10" swimtime="00:05:27.45" lane="5" heatid="10001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:11.95" />
                    <SPLIT distance="200" swimtime="00:02:36.48" />
                    <SPLIT distance="300" swimtime="00:04:02.20" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="496" eventid="18" swimtime="00:01:05.67" lane="4" heatid="18001" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="160" birthdate="2007-01-01" gender="M" lastname="Kühne" firstname="Gustav" license="0">
              <RESULTS>
                <RESULT resultid="498" eventid="9" status="DSQ" swimtime="00:00:59.18" lane="4" heatid="9005" comment="falsche Ausrüstung (Hose)" />
                <RESULT resultid="499" eventid="12" status="DSQ" swimtime="00:00:26.59" lane="1" heatid="12004" comment="falscher Start" />
                <RESULT resultid="500" eventid="14" swimtime="00:02:23.47" lane="3" heatid="14003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:09.81" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="161" birthdate="2008-01-01" gender="M" lastname="Steininger" firstname="Bruno" license="0">
              <RESULTS>
                <RESULT resultid="501" eventid="2" swimtime="00:00:20.35" lane="4" heatid="2002" />
                <RESULT resultid="502" eventid="14" swimtime="00:02:00.00" lane="3" heatid="14004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:56.13" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="503" eventid="17" swimtime="00:04:18.00" lane="8" heatid="17003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:01.27" />
                    <SPLIT distance="200" swimtime="00:02:09.47" />
                    <SPLIT distance="300" swimtime="00:03:17.04" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="504" eventid="19" swimtime="00:00:53.59" lane="3" heatid="19002" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="162" birthdate="2008-01-01" gender="F" lastname="Durcak" firstname="Clara" license="0">
              <RESULTS>
                <RESULT resultid="505" eventid="1" swimtime="00:00:28.17" lane="2" heatid="1002" />
                <RESULT resultid="506" eventid="8" swimtime="00:01:05.24" lane="2" heatid="8007" />
                <RESULT resultid="507" eventid="13" swimtime="00:02:24.87" lane="3" heatid="13006">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:08.46" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="508" eventid="18" swimtime="00:01:10.94" lane="8" heatid="18002" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="163" birthdate="2008-01-01" gender="F" lastname="Altenstein" firstname="Isabelle" license="0">
              <RESULTS>
                <RESULT resultid="509" eventid="1" swimtime="00:00:26.01" lane="7" heatid="1002" />
                <RESULT resultid="510" eventid="8" swimtime="00:01:00.80" lane="5" heatid="8007" />
                <RESULT resultid="511" eventid="11" swimtime="00:00:27.62" lane="2" heatid="11008" />
                <RESULT resultid="512" eventid="16" swimtime="00:04:52.55" lane="5" heatid="16003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:07.70" />
                    <SPLIT distance="200" swimtime="00:02:23.19" />
                    <SPLIT distance="300" swimtime="00:03:39.43" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="164" birthdate="2009-01-01" gender="F" lastname="Fabian" firstname="Ileen" license="0">
              <RESULTS>
                <RESULT resultid="513" eventid="8" swimtime="00:01:13.88" lane="6" heatid="8007" />
                <RESULT resultid="514" eventid="11" swimtime="00:00:29.28" lane="5" heatid="11007" />
                <RESULT resultid="515" eventid="13" swimtime="00:02:44.05" lane="8" heatid="13004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:15.66" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="516" eventid="18" swimtime="00:01:37.29" lane="3" heatid="18001" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="165" birthdate="2009-01-01" gender="F" lastname="Steininger" firstname="Magda" license="0">
              <RESULTS>
                <RESULT resultid="517" eventid="1" swimtime="00:00:24.47" lane="5" heatid="1002" />
                <RESULT resultid="518" eventid="11" swimtime="00:00:26.18" lane="4" heatid="11009" />
                <RESULT resultid="519" eventid="16" swimtime="00:04:55.47" lane="8" heatid="16004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:06.34" />
                    <SPLIT distance="200" swimtime="00:02:21.56" />
                    <SPLIT distance="300" swimtime="00:03:40.26" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="520" eventid="18" swimtime="00:01:03.03" lane="1" heatid="18002" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="166" birthdate="2012-01-01" gender="M" lastname="Gerbach" firstname="Linus" license="0">
              <RESULTS>
                <RESULT resultid="521" eventid="14" swimtime="00:03:02.67" lane="1" heatid="14002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:29.66" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="522" eventid="17" swimtime="00:06:07.14" lane="4" heatid="17001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:24.06" />
                    <SPLIT distance="200" swimtime="00:02:58.79" />
                    <SPLIT distance="300" swimtime="00:04:34.16" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="167" birthdate="2014-01-01" gender="F" lastname="Teufel" firstname="Sophia" license="0">
              <RESULTS>
                <RESULT resultid="523" eventid="5" swimtime="00:00:49.60" lane="5" heatid="5002" />
                <RESULT resultid="524" eventid="8" swimtime="00:01:37.29" lane="8" heatid="8003" />
                <RESULT resultid="525" eventid="11" status="DSQ" swimtime="00:00:43.68" lane="7" heatid="11003" comment="falscher Start" />
                <RESULT resultid="526" eventid="13" swimtime="00:03:30.08" lane="5" heatid="13002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:38.75" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY number="1" gender="F" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="477" eventid="20" swimtime="00:03:42.88" lane="2" heatid="20003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:52.81" />
                    <SPLIT distance="200" swimtime="00:01:51.79" />
                    <SPLIT distance="300" swimtime="00:02:51.75" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="152" number="1" />
                    <RELAYPOSITION athleteid="157" number="2" />
                    <RELAYPOSITION athleteid="165" number="3" />
                    <RELAYPOSITION athleteid="154" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" gender="M" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="488" eventid="21" status="EXH" swimtime="00:04:24.71" lane="2" heatid="21001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:51.69" />
                    <SPLIT distance="200" swimtime="00:02:01.77" />
                    <SPLIT distance="300" swimtime="00:03:25.69" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="161" number="1" />
                    <RELAYPOSITION athleteid="151" number="2" />
                    <RELAYPOSITION athleteid="166" number="3" />
                    <RELAYPOSITION athleteid="160" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" gender="F" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="497" eventid="20" swimtime="00:04:22.56" lane="4" heatid="20002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:02.19" />
                    <SPLIT distance="200" swimtime="00:02:15.83" />
                    <SPLIT distance="300" swimtime="00:03:22.76" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="158" number="1" />
                    <RELAYPOSITION athleteid="164" number="2" />
                    <RELAYPOSITION athleteid="162" number="3" />
                    <RELAYPOSITION athleteid="163" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB name="SSV Freiburg" nation="GER" region="33" code="0">
          <ATHLETES>
            <ATHLETE athleteid="14" birthdate="2000-01-01" gender="F" lastname="Köhn" firstname="Theresa" license="0">
              <RESULTS>
                <RESULT resultid="57" eventid="1" swimtime="00:00:20.61" lane="3" heatid="1006" />
                <RESULT resultid="52" eventid="8" swimtime="00:00:49.22" lane="5" heatid="8013" />
                <RESULT resultid="55" eventid="10" swimtime="00:03:54.09" lane="8" heatid="10003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:54.73" />
                    <SPLIT distance="200" swimtime="00:01:54.41" />
                    <SPLIT distance="300" swimtime="00:02:55.50" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="53" eventid="18" swimtime="00:00:47.55" lane="5" heatid="18004" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="15" birthdate="1998-01-01" gender="F" lastname="Köhn" firstname="Johanna" license="0">
              <RESULTS>
                <RESULT resultid="58" eventid="7" swimtime="00:08:21.08" lane="2" heatid="7004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:58.43" />
                    <SPLIT distance="200" swimtime="00:02:00.05" />
                    <SPLIT distance="300" swimtime="00:03:02.57" />
                    <SPLIT distance="400" swimtime="00:04:05.88" />
                    <SPLIT distance="500" swimtime="00:05:09.53" />
                    <SPLIT distance="600" swimtime="00:06:13.72" />
                    <SPLIT distance="700" swimtime="00:07:18.19" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="56" eventid="10" swimtime="00:03:50.79" lane="4" heatid="10002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:54.49" />
                    <SPLIT distance="200" swimtime="00:01:52.59" />
                    <SPLIT distance="300" swimtime="00:02:52.15" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="54" eventid="16" swimtime="00:04:08.11" lane="8" heatid="16008">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:58.92" />
                    <SPLIT distance="200" swimtime="00:02:01.98" />
                    <SPLIT distance="300" swimtime="00:03:05.56" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="Tauchclub Heilbronn" nation="GER" region="32" code="0">
          <ATHLETES>
            <ATHLETE athleteid="16" birthdate="2004-01-01" gender="F" lastname="Ruedel" firstname="Leona" license="0">
              <RESULTS>
                <RESULT resultid="91" eventid="1" swimtime="00:00:20.65" lane="4" heatid="1005" />
                <RESULT resultid="59" eventid="8" swimtime="00:00:48.78" lane="7" heatid="8013" />
                <RESULT resultid="101" eventid="11" swimtime="00:00:22.48" lane="3" heatid="11013" />
                <RESULT resultid="75" eventid="13" swimtime="00:01:51.48" lane="6" heatid="13009">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:54.45" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="70" eventid="18" swimtime="00:00:52.77" lane="1" heatid="18004" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="17" birthdate="2004-01-01" gender="F" lastname="Phillipp" firstname="Beeke Alea" license="0">
              <RESULTS>
                <RESULT resultid="92" eventid="1" swimtime="00:00:20.86" lane="3" heatid="1005" />
                <RESULT resultid="60" eventid="8" swimtime="00:00:51.77" lane="1" heatid="8013" />
                <RESULT resultid="102" eventid="11" swimtime="00:00:22.86" lane="7" heatid="11013" />
                <RESULT resultid="74" eventid="13" swimtime="00:01:58.02" lane="8" heatid="13010">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:54.92" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="69" eventid="18" swimtime="00:00:50.12" lane="2" heatid="18004" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="18" birthdate="2008-01-01" gender="F" lastname="Seidel" firstname="Esther-Sophie" license="0">
              <RESULTS>
                <RESULT resultid="93" eventid="1" swimtime="00:00:22.27" lane="7" heatid="1004" />
                <RESULT resultid="61" eventid="8" swimtime="00:00:56.40" lane="5" heatid="8011" />
                <RESULT resultid="104" eventid="11" swimtime="00:00:24.18" lane="8" heatid="11012" />
                <RESULT resultid="78" eventid="13" swimtime="00:02:09.85" lane="2" heatid="13007">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:04.22" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="85" eventid="16" swimtime="00:04:42.24" lane="7" heatid="16004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:05.65" />
                    <SPLIT distance="200" swimtime="00:02:20.05" />
                    <SPLIT distance="300" swimtime="00:03:32.41" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="19" birthdate="2009-01-01" gender="F" lastname="Hölzer" firstname="Elisa" license="0">
              <RESULTS>
                <RESULT resultid="94" eventid="1" swimtime="00:00:22.81" lane="1" heatid="1004" />
                <RESULT resultid="62" eventid="8" swimtime="00:00:54.15" lane="2" heatid="8011" />
                <RESULT resultid="103" eventid="11" swimtime="00:00:24.19" lane="3" heatid="11012" />
                <RESULT resultid="76" eventid="13" swimtime="00:02:02.83" lane="7" heatid="13008">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:57.65" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="83" eventid="16" swimtime="00:04:28.25" lane="3" heatid="16005">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:01.81" />
                    <SPLIT distance="200" swimtime="00:02:10.53" />
                    <SPLIT distance="300" swimtime="00:03:21.31" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="20" birthdate="2009-01-01" gender="F" lastname="Rettig" firstname="Sina" license="0">
              <RESULTS>
                <RESULT resultid="96" eventid="1" swimtime="00:00:24.41" lane="8" heatid="1003" />
                <RESULT resultid="63" eventid="8" swimtime="00:01:00.00" lane="7" heatid="8010" />
                <RESULT resultid="105" eventid="11" swimtime="00:00:25.77" lane="2" heatid="11010" />
                <RESULT resultid="79" eventid="13" swimtime="00:02:19.79" lane="4" heatid="13006">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:05.74" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="86" eventid="16" swimtime="00:05:05.78" lane="4" heatid="16003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:09.04" />
                    <SPLIT distance="200" swimtime="00:02:28.32" />
                    <SPLIT distance="300" swimtime="00:03:49.71" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="21" birthdate="2008-01-01" gender="F" lastname="Grimm" firstname="Hannah" license="0">
              <RESULTS>
                <RESULT resultid="95" eventid="1" swimtime="00:00:24.19" lane="5" heatid="1003" />
                <RESULT resultid="64" eventid="8" swimtime="00:00:57.18" lane="5" heatid="8009" />
                <RESULT resultid="106" eventid="11" swimtime="00:00:25.34" lane="7" heatid="11010" />
                <RESULT resultid="77" eventid="13" swimtime="00:02:10.82" lane="3" heatid="13007">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:02.29" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="84" eventid="16" swimtime="00:04:41.88" lane="4" heatid="16004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:05.82" />
                    <SPLIT distance="200" swimtime="00:02:19.01" />
                    <SPLIT distance="300" swimtime="00:03:34.20" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="22" birthdate="2003-01-01" gender="M" lastname="Fabriz" firstname="Tobias" license="0">
              <RESULTS>
                <RESULT resultid="97" eventid="2" swimtime="00:00:17.96" lane="1" heatid="2006" />
                <RESULT resultid="65" eventid="9" swimtime="00:00:46.01" lane="7" heatid="9009" />
                <RESULT resultid="107" eventid="12" status="DNS" swimtime="00:00:00.00" lane="3" heatid="12008" />
                <RESULT resultid="71" eventid="19" status="DNS" swimtime="00:00:00.00" lane="1" heatid="19004" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="23" birthdate="2007-01-01" gender="M" lastname="Bilicz" firstname="Benedikt" license="0">
              <RESULTS>
                <RESULT resultid="98" eventid="2" swimtime="00:00:19.27" lane="5" heatid="2004" />
                <RESULT resultid="66" eventid="9" status="DSQ" swimtime="00:00:48.91" lane="2" heatid="9008" comment="15m nach Start übertaucht" />
                <RESULT resultid="108" eventid="12" swimtime="00:00:21.88" lane="6" heatid="12007" />
                <RESULT resultid="80" eventid="14" swimtime="00:01:52.96" lane="6" heatid="14005">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:53.71" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="72" eventid="19" swimtime="00:00:49.37" lane="8" heatid="19003" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="24" birthdate="2002-01-01" gender="M" lastname="Bauer" firstname="Sebastian" license="0">
              <RESULTS>
                <RESULT resultid="99" eventid="2" swimtime="00:00:19.94" lane="8" heatid="2004" />
                <RESULT resultid="67" eventid="9" swimtime="00:00:51.89" lane="5" heatid="9007" />
                <RESULT resultid="109" eventid="12" swimtime="00:00:23.59" lane="8" heatid="12007" />
                <RESULT resultid="87" eventid="17" swimtime="00:04:19.65" lane="8" heatid="17004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:57.45" />
                    <SPLIT distance="200" swimtime="00:02:02.61" />
                    <SPLIT distance="300" swimtime="00:03:11.42" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="25" birthdate="2011-01-01" gender="M" lastname="Korb" firstname="Elias" license="0">
              <RESULTS>
                <RESULT resultid="111" eventid="4" swimtime="00:00:25.63" lane="5" heatid="4002" />
                <RESULT resultid="68" eventid="9" swimtime="00:00:58.46" lane="7" heatid="9006" />
                <RESULT resultid="110" eventid="12" swimtime="00:00:26.23" lane="6" heatid="12005" />
                <RESULT resultid="82" eventid="14" swimtime="00:02:08.43" lane="2" heatid="14004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:02.82" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="73" eventid="19" swimtime="00:00:58.97" lane="7" heatid="19002" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="26" birthdate="2004-01-01" gender="M" lastname="Rist" firstname="Marc" license="0">
              <RESULTS>
                <RESULT resultid="100" eventid="2" swimtime="00:00:22.50" lane="8" heatid="2003" />
                <RESULT resultid="112" eventid="7" swimtime="00:09:05.09" lane="6" heatid="7002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:59.31" />
                    <SPLIT distance="200" swimtime="00:02:07.59" />
                    <SPLIT distance="300" swimtime="00:03:17.43" />
                    <SPLIT distance="400" swimtime="00:04:27.54" />
                    <SPLIT distance="500" swimtime="00:05:39.25" />
                    <SPLIT distance="600" swimtime="00:06:50.60" />
                    <SPLIT distance="700" swimtime="00:08:00.35" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="81" eventid="14" swimtime="00:01:54.54" lane="2" heatid="14005">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:55.63" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="88" eventid="17" swimtime="00:04:16.77" lane="6" heatid="17003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:58.69" />
                    <SPLIT distance="200" swimtime="00:02:05.32" />
                    <SPLIT distance="300" swimtime="00:03:13.42" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY number="1" gender="F" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="89" eventid="20" swimtime="00:03:49.65" lane="5" heatid="20003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:53.42" />
                    <SPLIT distance="200" swimtime="00:01:51.70" />
                    <SPLIT distance="300" swimtime="00:02:55.06" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="18" number="1" />
                    <RELAYPOSITION athleteid="21" number="2" />
                    <RELAYPOSITION athleteid="20" number="3" />
                    <RELAYPOSITION athleteid="19" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" gender="M" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="90" eventid="21" swimtime="00:03:33.15" lane="6" heatid="21002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:51.82" />
                    <SPLIT distance="200" swimtime="00:01:45.43" />
                    <SPLIT distance="300" swimtime="00:02:34.35" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="26" number="1" />
                    <RELAYPOSITION athleteid="24" number="2" />
                    <RELAYPOSITION athleteid="23" number="3" />
                    <RELAYPOSITION athleteid="25" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB name="Tauchclub NEMO Plauen e.V." nation="GER" region="20" code="0">
          <ATHLETES>
            <ATHLETE athleteid="37" birthdate="2012-01-01" gender="F" lastname="Troppschuh" firstname="Lotte" license="0">
              <RESULTS>
                <RESULT resultid="134" eventid="8" swimtime="00:00:54.07" lane="7" heatid="8011" />
                <RESULT resultid="139" eventid="11" swimtime="00:00:23.99" lane="5" heatid="11012" />
                <RESULT resultid="136" eventid="16" swimtime="00:04:52.15" lane="8" heatid="16005">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:03.81" />
                    <SPLIT distance="200" swimtime="00:02:20.28" />
                    <SPLIT distance="300" swimtime="00:03:38.67" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="38" birthdate="2009-01-01" gender="F" lastname="Troppschuh" firstname="Hannah" license="0">
              <RESULTS>
                <RESULT resultid="137" eventid="1" swimtime="00:00:18.78" lane="2" heatid="1006" />
                <RESULT resultid="138" eventid="11" swimtime="00:00:21.86" lane="8" heatid="11014" />
                <RESULT resultid="135" eventid="18" swimtime="00:00:43.93" lane="1" heatid="18005" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="Tauchsportclub Erfurt e.V." nation="GER" region="35" code="0">
          <ATHLETES>
            <ATHLETE athleteid="220" birthdate="2011-01-01" gender="F" lastname="Döll" firstname="Katharina Martha" license="0">
              <RESULTS>
                <RESULT resultid="691" eventid="8" swimtime="00:01:20.07" lane="5" heatid="8001" />
                <RESULT resultid="780" eventid="11" swimtime="00:00:34.77" lane="6" heatid="11001" />
                <RESULT resultid="729" eventid="13" swimtime="00:03:06.87" lane="5" heatid="13001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:26.19" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="221" birthdate="2003-01-01" gender="F" lastname="Thomas" firstname="Nina" license="0">
              <RESULTS>
                <RESULT resultid="764" eventid="1" swimtime="00:00:22.47" lane="4" heatid="1004" />
                <RESULT resultid="692" eventid="8" swimtime="00:00:52.31" lane="1" heatid="8012" />
                <RESULT resultid="730" eventid="13" swimtime="00:02:01.34" lane="7" heatid="13009">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:57.98" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="747" eventid="16" swimtime="00:04:27.58" lane="7" heatid="16006">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:02.65" />
                    <SPLIT distance="200" swimtime="00:02:12.27" />
                    <SPLIT distance="300" swimtime="00:03:21.11" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="222" birthdate="2010-01-01" gender="F" lastname="Abe" firstname="Adina" license="0">
              <RESULTS>
                <RESULT resultid="809" eventid="3" swimtime="00:00:25.03" lane="4" heatid="3001" />
                <RESULT resultid="693" eventid="8" swimtime="00:00:55.09" lane="6" heatid="8011" />
                <RESULT resultid="782" eventid="11" swimtime="00:00:25.30" lane="4" heatid="11011" />
                <RESULT resultid="731" eventid="13" swimtime="00:02:03.84" lane="2" heatid="13008">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:00.05" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="720" eventid="18" swimtime="00:00:57.55" lane="1" heatid="18003" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="223" birthdate="2009-01-01" gender="F" lastname="Zitzmann" firstname="Annalena" license="0">
              <RESULTS>
                <RESULT resultid="767" eventid="1" swimtime="00:00:23.84" lane="6" heatid="1002" />
                <RESULT resultid="694" eventid="8" swimtime="00:00:55.99" lane="1" heatid="8011" />
                <RESULT resultid="783" eventid="11" swimtime="00:00:24.88" lane="5" heatid="11011" />
                <RESULT resultid="732" eventid="13" swimtime="00:02:07.20" lane="4" heatid="13007">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:01.16" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="721" eventid="18" swimtime="00:00:57.48" lane="8" heatid="18003" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="224" birthdate="2004-01-01" gender="F" lastname="Möller" firstname="Amelie" license="0">
              <RESULTS>
                <RESULT resultid="695" eventid="8" status="DSQ" swimtime="00:00:58.10" lane="8" heatid="8011" comment="falscher Start" />
                <RESULT resultid="784" eventid="11" swimtime="00:00:25.91" lane="8" heatid="11011" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="225" birthdate="1979-01-01" gender="F" lastname="Leipold" firstname="Steffi" license="0">
              <RESULTS>
                <RESULT resultid="696" eventid="8" swimtime="00:00:59.01" lane="3" heatid="8009" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="226" birthdate="1982-01-01" gender="F" lastname="Zitzmann" firstname="Ulrike" license="0">
              <RESULTS>
                <RESULT resultid="697" eventid="8" swimtime="00:01:03.74" lane="5" heatid="8008" />
                <RESULT resultid="788" eventid="11" swimtime="00:00:28.89" lane="8" heatid="11008" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="227" birthdate="2006-01-01" gender="F" lastname="Heinitz" firstname="Leonor" license="0">
              <RESULTS>
                <RESULT resultid="766" eventid="1" swimtime="00:00:22.29" lane="3" heatid="1002" />
                <RESULT resultid="698" eventid="8" swimtime="00:00:55.78" lane="3" heatid="8008" />
                <RESULT resultid="785" eventid="11" swimtime="00:00:25.36" lane="6" heatid="11009" />
                <RESULT resultid="733" eventid="13" swimtime="00:02:04.29" lane="6" heatid="13007">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:58.06" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="722" eventid="18" swimtime="00:00:55.77" lane="6" heatid="18002" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="228" birthdate="2007-01-01" gender="F" lastname="Zieger" firstname="Emilie" license="0">
              <RESULTS>
                <RESULT resultid="699" eventid="8" swimtime="00:01:07.05" lane="2" heatid="8008" />
                <RESULT resultid="787" eventid="11" swimtime="00:00:28.86" lane="7" heatid="11008" />
                <RESULT resultid="735" eventid="13" swimtime="00:02:22.67" lane="2" heatid="13006">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:07.18" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="229" birthdate="2009-01-01" gender="F" lastname="Henkel" firstname="Friederike" license="0">
              <RESULTS>
                <RESULT resultid="700" eventid="8" status="DNS" swimtime="00:00:00.00" lane="7" heatid="8008" />
                <RESULT resultid="786" eventid="11" status="DNS" swimtime="00:00:00.00" lane="8" heatid="11009" />
                <RESULT resultid="734" eventid="13" status="DNS" swimtime="00:00:00.00" lane="8" heatid="13007" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="230" birthdate="2009-01-01" gender="F" lastname="Blumenstein" firstname="Martha" license="0">
              <RESULTS>
                <RESULT resultid="768" eventid="1" swimtime="00:00:27.42" lane="1" heatid="1002" />
                <RESULT resultid="701" eventid="8" swimtime="00:00:59.33" lane="1" heatid="8008" />
                <RESULT resultid="748" eventid="16" swimtime="00:04:44.87" lane="6" heatid="16004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:05.92" />
                    <SPLIT distance="200" swimtime="00:02:20.26" />
                    <SPLIT distance="300" swimtime="00:03:34.49" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="728" eventid="22" swimtime="00:19:20.32" lane="3" heatid="22001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:08.24" />
                    <SPLIT distance="200" swimtime="00:02:25.56" />
                    <SPLIT distance="300" swimtime="00:03:43.11" />
                    <SPLIT distance="400" swimtime="00:05:01.60" />
                    <SPLIT distance="500" swimtime="00:06:19.39" />
                    <SPLIT distance="600" swimtime="00:07:37.87" />
                    <SPLIT distance="700" swimtime="00:08:55.80" />
                    <SPLIT distance="800" swimtime="00:10:14.79" />
                    <SPLIT distance="900" swimtime="00:11:33.95" />
                    <SPLIT distance="1000" swimtime="00:12:53.91" />
                    <SPLIT distance="1100" swimtime="00:14:13.17" />
                    <SPLIT distance="1200" swimtime="00:15:32.54" />
                    <SPLIT distance="1300" swimtime="00:16:51.16" />
                    <SPLIT distance="1400" swimtime="00:18:08.27" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="231" birthdate="2011-01-01" gender="F" lastname="Behrmann" firstname="Fine Erna" license="0">
              <RESULTS>
                <RESULT resultid="702" eventid="8" swimtime="00:01:06.42" lane="3" heatid="8007" />
                <RESULT resultid="789" eventid="11" swimtime="00:00:29.45" lane="6" heatid="11007" />
                <RESULT resultid="736" eventid="13" swimtime="00:02:38.91" lane="6" heatid="13005">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:13.63" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="232" birthdate="1968-01-01" gender="F" lastname="König" firstname="Sabine" license="0">
              <RESULTS>
                <RESULT resultid="703" eventid="8" swimtime="00:01:13.35" lane="4" heatid="8006" />
                <RESULT resultid="790" eventid="11" swimtime="00:00:32.56" lane="4" heatid="11006" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="233" birthdate="2012-01-01" gender="F" lastname="Blumenstein" firstname="Liese" license="0">
              <RESULTS>
                <RESULT resultid="776" eventid="5" swimtime="00:00:35.29" lane="1" heatid="5003" />
                <RESULT resultid="704" eventid="8" swimtime="00:01:12.97" lane="1" heatid="8006" />
                <RESULT resultid="793" eventid="11" swimtime="00:00:36.23" lane="5" heatid="11004" />
                <RESULT resultid="737" eventid="13" swimtime="00:02:41.85" lane="4" heatid="13004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:18.88" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="749" eventid="16" swimtime="00:05:43.64" lane="7" heatid="16003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:20.61" />
                    <SPLIT distance="200" swimtime="00:02:51.71" />
                    <SPLIT distance="300" swimtime="00:04:21.84" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="234" birthdate="2012-01-01" gender="F" lastname="Schulze" firstname="Paula" license="0">
              <RESULTS>
                <RESULT resultid="777" eventid="5" status="DSQ" swimtime="00:00:32.20" lane="4" heatid="5002" comment="falscher Stil über gesamte Strecke" />
                <RESULT resultid="705" eventid="8" swimtime="00:01:15.47" lane="5" heatid="8005" />
                <RESULT resultid="792" eventid="11" swimtime="00:00:32.58" lane="5" heatid="11005" />
                <RESULT resultid="738" eventid="13" swimtime="00:02:52.83" lane="6" heatid="13003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:23.13" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="751" eventid="16" status="DSQ" swimtime="00:00:00.00" lane="6" heatid="16002" comment="aufgegeben nach 250m">
                  <SPLITS>
                    <SPLIT distance="200" swimtime="00:01:33.59" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="235" birthdate="2010-01-01" gender="F" lastname="Hartung" firstname="Antonia" license="0">
              <RESULTS>
                <RESULT resultid="706" eventid="8" swimtime="00:01:24.30" lane="7" heatid="8005" />
                <RESULT resultid="791" eventid="11" swimtime="00:00:34.84" lane="3" heatid="11006" />
                <RESULT resultid="750" eventid="16" swimtime="00:06:38.70" lane="3" heatid="16002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:33.09" />
                    <SPLIT distance="200" swimtime="00:03:18.76" />
                    <SPLIT distance="300" swimtime="00:05:04.37" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="236" birthdate="2012-01-01" gender="F" lastname="Dallgas" firstname="Tia" license="0">
              <RESULTS>
                <RESULT resultid="775" eventid="5" swimtime="00:00:40.63" lane="2" heatid="5001" />
                <RESULT resultid="707" eventid="8" swimtime="00:01:27.29" lane="4" heatid="8002" />
                <RESULT resultid="794" eventid="11" swimtime="00:00:32.08" lane="1" heatid="11004" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="237" birthdate="2006-01-01" gender="M" lastname="Leipold" firstname="Marek" license="0">
              <RESULTS>
                <RESULT resultid="769" eventid="2" swimtime="00:00:15.79" lane="5" heatid="2006" />
                <RESULT resultid="708" eventid="9" swimtime="00:00:37.70" lane="5" heatid="9010" />
                <RESULT resultid="796" eventid="12" swimtime="00:00:16.92" lane="4" heatid="12009" />
                <RESULT resultid="724" eventid="19" swimtime="00:00:36.05" lane="3" heatid="19004" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="238" birthdate="1970-01-01" gender="M" lastname="Timpel" firstname="Heiko" license="0">
              <RESULTS>
                <RESULT resultid="770" eventid="2" swimtime="00:00:20.26" lane="1" heatid="2004" />
                <RESULT resultid="709" eventid="9" swimtime="00:00:49.75" lane="8" heatid="9008" />
                <RESULT resultid="797" eventid="12" swimtime="00:00:23.16" lane="4" heatid="12006" />
                <RESULT resultid="725" eventid="19" swimtime="00:00:45.41" lane="3" heatid="19003" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="239" birthdate="2008-01-01" gender="M" lastname="Hannemann" firstname="Fynn" license="0">
              <RESULTS>
                <RESULT resultid="771" eventid="2" swimtime="00:00:21.98" lane="5" heatid="2003" />
                <RESULT resultid="710" eventid="9" swimtime="00:00:51.96" lane="6" heatid="9007" />
                <RESULT resultid="798" eventid="12" swimtime="00:00:23.47" lane="3" heatid="12006" />
                <RESULT resultid="739" eventid="14" swimtime="00:02:08.40" lane="8" heatid="14005">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:02.11" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="727" eventid="19" swimtime="00:00:55.99" lane="2" heatid="19002" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="240" birthdate="2010-01-01" gender="M" lastname="Leipold" firstname="Jakob" license="0">
              <RESULTS>
                <RESULT resultid="812" eventid="4" swimtime="00:00:24.37" lane="4" heatid="4002" />
                <RESULT resultid="711" eventid="9" swimtime="00:00:56.42" lane="5" heatid="9006" />
                <RESULT resultid="799" eventid="12" swimtime="00:00:26.57" lane="7" heatid="12006" />
                <RESULT resultid="740" eventid="14" swimtime="00:02:08.04" lane="5" heatid="14004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:01.98" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="726" eventid="19" swimtime="00:00:59.30" lane="5" heatid="19002" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="241" birthdate="1978-01-01" gender="M" lastname="Hannemann" firstname="Ronny" license="0">
              <RESULTS>
                <RESULT resultid="772" eventid="2" swimtime="00:00:24.24" lane="3" heatid="2002" />
                <RESULT resultid="712" eventid="9" swimtime="00:00:56.32" lane="2" heatid="9006" />
                <RESULT resultid="800" eventid="12" swimtime="00:00:26.03" lane="5" heatid="12005" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="242" birthdate="2010-01-01" gender="M" lastname="Hochstein" firstname="Jean Paul" license="0">
              <RESULTS>
                <RESULT resultid="810" eventid="4" swimtime="00:00:30.95" lane="4" heatid="4001" />
                <RESULT resultid="713" eventid="9" swimtime="00:01:00.94" lane="3" heatid="9005" />
                <RESULT resultid="802" eventid="12" swimtime="00:00:26.96" lane="5" heatid="12004" />
                <RESULT resultid="742" eventid="14" swimtime="00:02:18.79" lane="5" heatid="14003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:07.20" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="753" eventid="17" swimtime="00:05:15.99" lane="6" heatid="17002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:15.81" />
                    <SPLIT distance="200" swimtime="00:02:40.63" />
                    <SPLIT distance="300" swimtime="00:04:04.54" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="243" birthdate="1971-01-01" gender="M" lastname="Schmidt" firstname="Alexander" license="0">
              <RESULTS>
                <RESULT resultid="773" eventid="2" swimtime="00:00:29.72" lane="4" heatid="2001" />
                <RESULT resultid="714" eventid="9" swimtime="00:01:02.68" lane="6" heatid="9005" />
                <RESULT resultid="801" eventid="12" swimtime="00:00:27.53" lane="8" heatid="12005" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="244" birthdate="2010-01-01" gender="M" lastname="Hochstein" firstname="Maddox Lee" license="0">
              <RESULTS>
                <RESULT resultid="811" eventid="4" swimtime="00:00:26.99" lane="7" heatid="4002" />
                <RESULT resultid="715" eventid="9" swimtime="00:01:02.09" lane="1" heatid="9005" />
                <RESULT resultid="803" eventid="12" swimtime="00:00:26.45" lane="3" heatid="12004" />
                <RESULT resultid="741" eventid="14" swimtime="00:02:19.72" lane="8" heatid="14004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:07.86" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="752" eventid="17" swimtime="00:05:04.60" lane="3" heatid="17002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:09.78" />
                    <SPLIT distance="200" swimtime="00:02:28.79" />
                    <SPLIT distance="300" swimtime="00:03:50.02" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="245" birthdate="2010-01-01" gender="M" lastname="Blumenstein" firstname="Einar" license="0">
              <RESULTS>
                <RESULT resultid="716" eventid="9" status="DSQ" swimtime="00:01:13.61" lane="1" heatid="9004" comment="falscher Start" />
                <RESULT resultid="805" eventid="12" swimtime="00:00:30.57" lane="5" heatid="12003" />
                <RESULT resultid="744" eventid="14" status="DSQ" swimtime="00:00:00.00" lane="8" heatid="14003" comment="aufgegeben nach 150m">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:10.86" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="246" birthdate="2010-01-01" gender="M" lastname="Schmidt" firstname="Jakob" license="0">
              <RESULTS>
                <RESULT resultid="717" eventid="9" swimtime="00:01:15.72" lane="2" heatid="9003" />
                <RESULT resultid="806" eventid="12" swimtime="00:00:34.68" lane="8" heatid="12003" />
                <RESULT resultid="745" eventid="14" swimtime="00:02:55.48" lane="4" heatid="14001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:23.72" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="249" birthdate="2009-01-01" gender="M" lastname="Artschwager" firstname="Gustaf" license="0">
              <RESULTS>
                <RESULT resultid="814" eventid="7" swimtime="00:10:50.75" lane="3" heatid="7001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:11.18" />
                    <SPLIT distance="200" swimtime="00:02:34.13" />
                    <SPLIT distance="300" swimtime="00:03:59.43" />
                    <SPLIT distance="400" swimtime="00:05:25.30" />
                    <SPLIT distance="500" swimtime="00:06:51.15" />
                    <SPLIT distance="600" swimtime="00:08:14.19" />
                    <SPLIT distance="700" swimtime="00:09:36.86" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="804" eventid="12" swimtime="00:00:27.25" lane="7" heatid="12004" />
                <RESULT resultid="743" eventid="14" swimtime="00:02:18.19" lane="7" heatid="14003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:07.18" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="723" eventid="19" swimtime="00:01:13.51" lane="6" heatid="19001" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="258" birthdate="2009-01-01" gender="F" lastname="Darzhaniia" firstname="Alisa" license="0">
              <RESULTS>
                <RESULT resultid="765" eventid="1" swimtime="00:00:20.06" lane="3" heatid="1004" />
                <RESULT resultid="813" eventid="7" swimtime="00:08:45.02" lane="6" heatid="7003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:58.22" />
                    <SPLIT distance="200" swimtime="00:02:03.36" />
                    <SPLIT distance="300" swimtime="00:03:10.64" />
                    <SPLIT distance="400" swimtime="00:04:18.91" />
                    <SPLIT distance="500" swimtime="00:05:28.78" />
                    <SPLIT distance="600" swimtime="00:06:37.54" />
                    <SPLIT distance="700" swimtime="00:07:44.28" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="781" eventid="11" swimtime="00:00:22.11" lane="5" heatid="11013" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="259" birthdate="2013-01-01" gender="F" lastname="Medola" firstname="Anna" license="0">
              <RESULTS>
                <RESULT resultid="774" eventid="5" swimtime="00:00:46.09" lane="6" heatid="5001" />
                <RESULT resultid="795" eventid="11" status="DSQ" swimtime="00:00:39.13" lane="3" heatid="11002" comment="falscher Start" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="260" birthdate="1976-01-01" gender="F" lastname="Zieger" firstname="Katrin" license="0" />
            <ATHLETE athleteid="261" birthdate="1977-01-01" gender="F" lastname="Blumenstein" firstname="Sandra" license="0" />
            <ATHLETE athleteid="262" birthdate="1979-01-01" gender="F" lastname="Möller" firstname="Susanne" license="0" />
            <ATHLETE athleteid="311" birthdate="2009-01-01" gender="F" lastname="Naupold" firstname="Celina" license="0" />
          </ATHLETES>
          <RELAYS>
            <RELAY number="1" gender="F" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="754" eventid="20" swimtime="00:03:36.97" lane="8" heatid="20003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:49.47" />
                    <SPLIT distance="200" swimtime="00:01:45.03" />
                    <SPLIT distance="300" swimtime="00:02:40.87" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="258" number="1" />
                    <RELAYPOSITION athleteid="222" number="2" />
                    <RELAYPOSITION athleteid="223" number="3" />
                    <RELAYPOSITION athleteid="227" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="2" gender="F" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="755" eventid="20" status="EXH" swimtime="00:04:17.57" lane="5" heatid="20002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:12.14" />
                    <SPLIT distance="200" swimtime="00:02:09.47" />
                    <SPLIT distance="300" swimtime="00:03:11.94" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="228" number="1" />
                    <RELAYPOSITION athleteid="311" number="2" />
                    <RELAYPOSITION athleteid="230" number="3" />
                    <RELAYPOSITION athleteid="231" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="3" gender="F" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="756" eventid="20" swimtime="00:05:12.33" lane="4" heatid="20001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:14.24" />
                    <SPLIT distance="200" swimtime="00:02:30.62" />
                    <SPLIT distance="300" swimtime="00:03:52.19" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="233" number="1" />
                    <RELAYPOSITION athleteid="234" number="2" />
                    <RELAYPOSITION athleteid="220" number="3" />
                    <RELAYPOSITION athleteid="235" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" gender="X" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="761" eventid="15" swimtime="00:01:48.35" lane="4" heatid="15002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:50.13" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="243" number="1" />
                    <RELAYPOSITION athleteid="238" number="2" />
                    <RELAYPOSITION athleteid="225" number="3" />
                    <RELAYPOSITION athleteid="232" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" gender="X" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="762" eventid="15" swimtime="00:01:56.72" lane="3" heatid="15002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:56.51" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="241" number="1" />
                    <RELAYPOSITION athleteid="260" number="2" />
                    <RELAYPOSITION athleteid="262" number="3" />
                    <RELAYPOSITION athleteid="226" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" gender="M" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="759" eventid="21" swimtime="00:03:35.44" lane="7" heatid="21002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:40.83" />
                    <SPLIT distance="200" swimtime="00:01:36.48" />
                    <SPLIT distance="300" swimtime="00:02:33.76" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="237" number="1" />
                    <RELAYPOSITION athleteid="239" number="2" />
                    <RELAYPOSITION athleteid="240" number="3" />
                    <RELAYPOSITION athleteid="242" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="2" gender="M" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="760" eventid="21" swimtime="00:04:32.73" lane="7" heatid="21001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:03.22" />
                    <SPLIT distance="200" swimtime="00:02:05.93" />
                    <SPLIT distance="300" swimtime="00:03:14.76" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="249" number="1" />
                    <RELAYPOSITION athleteid="244" number="2" />
                    <RELAYPOSITION athleteid="245" number="3" />
                    <RELAYPOSITION athleteid="246" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" gender="X" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="763" eventid="15" swimtime="00:02:17.35" lane="3" heatid="15001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:05.47" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="234" number="1" />
                    <RELAYPOSITION athleteid="236" number="2" />
                    <RELAYPOSITION athleteid="259" number="3" />
                    <RELAYPOSITION athleteid="233" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" gender="X" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="815" eventid="21" swimtime="00:04:22.46" lane="3" heatid="21001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:06.02" />
                    <SPLIT distance="200" swimtime="00:02:11.72" />
                    <SPLIT distance="300" swimtime="00:03:26.36" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="260" number="1" />
                    <RELAYPOSITION athleteid="226" number="2" />
                    <RELAYPOSITION athleteid="262" number="3" />
                    <RELAYPOSITION athleteid="241" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" gender="X" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="816" eventid="21" swimtime="00:04:08.33" lane="4" heatid="21001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:59.70" />
                    <SPLIT distance="200" swimtime="00:02:01.05" />
                    <SPLIT distance="300" swimtime="00:03:17.25" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="225" number="1" />
                    <RELAYPOSITION athleteid="243" number="2" />
                    <RELAYPOSITION athleteid="232" number="3" />
                    <RELAYPOSITION athleteid="238" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB name="TC Chemie Greiz e.V." nation="GER" region="35" code="0">
          <ATHLETES>
            <ATHLETE athleteid="177" birthdate="1974-01-01" gender="M" lastname="Kühn" firstname="Ronald" license="0">
              <RESULTS>
                <RESULT resultid="555" eventid="2" swimtime="00:00:21.92" lane="7" heatid="2003" />
                <RESULT resultid="556" eventid="9" swimtime="00:00:56.07" lane="4" heatid="9006" />
                <RESULT resultid="557" eventid="12" swimtime="00:00:25.17" lane="1" heatid="12006" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="179" birthdate="2005-01-01" gender="F" lastname="Kupka" firstname="Miriam" license="0">
              <RESULTS>
                <RESULT resultid="563" eventid="1" swimtime="00:00:19.12" lane="7" heatid="1006" />
                <RESULT resultid="564" eventid="8" swimtime="00:00:46.32" lane="4" heatid="8013" />
                <RESULT resultid="565" eventid="11" swimtime="00:00:20.65" lane="4" heatid="11013" />
                <RESULT resultid="566" eventid="13" swimtime="00:01:48.48" lane="1" heatid="13011">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:51.23" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="567" eventid="16" swimtime="00:04:06.25" lane="3" heatid="16007">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:56.91" />
                    <SPLIT distance="200" swimtime="00:02:00.25" />
                    <SPLIT distance="300" swimtime="00:03:05.24" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="181" birthdate="2006-01-01" gender="F" lastname="Frauenfelder" firstname="Anneliese" license="0">
              <RESULTS>
                <RESULT resultid="569" eventid="1" swimtime="00:00:20.42" lane="8" heatid="1006" />
                <RESULT resultid="570" eventid="8" swimtime="00:00:49.57" lane="8" heatid="8013" />
                <RESULT resultid="571" eventid="10" swimtime="00:04:23.54" lane="3" heatid="10002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:57.74" />
                    <SPLIT distance="200" swimtime="00:02:03.67" />
                    <SPLIT distance="300" swimtime="00:03:13.69" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="572" eventid="18" swimtime="00:00:46.82" lane="8" heatid="18005" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="183" birthdate="2008-01-01" gender="M" lastname="Lose" firstname="Fabian" license="0">
              <RESULTS>
                <RESULT resultid="577" eventid="9" swimtime="00:00:59.07" lane="2" heatid="9005" />
                <RESULT resultid="578" eventid="12" swimtime="00:00:27.19" lane="6" heatid="12004" />
                <RESULT resultid="579" eventid="14" status="DSQ" swimtime="00:02:16.71" lane="6" heatid="14003" comment="falscher Start">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:07.85" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="580" eventid="19" swimtime="00:01:07.30" lane="6" heatid="19002" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="184" birthdate="2008-01-01" gender="M" lastname="Robenz" firstname="Jean Robin" license="0">
              <RESULTS>
                <RESULT resultid="581" eventid="2" swimtime="00:00:27.37" lane="7" heatid="2001" />
                <RESULT resultid="582" eventid="9" swimtime="00:01:01.47" lane="3" heatid="9004" />
                <RESULT resultid="583" eventid="12" swimtime="00:00:27.05" lane="7" heatid="12002" />
                <RESULT resultid="584" eventid="14" swimtime="00:02:16.32" lane="1" heatid="14003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:04.37" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="585" eventid="19" swimtime="00:01:05.67" lane="5" heatid="19001" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="185" birthdate="2008-01-01" gender="M" lastname="Berger" firstname="Louis" license="0">
              <RESULTS>
                <RESULT resultid="586" eventid="9" swimtime="00:00:44.20" lane="3" heatid="9009" />
                <RESULT resultid="587" eventid="12" swimtime="00:00:19.85" lane="8" heatid="12009" />
                <RESULT resultid="588" eventid="14" swimtime="00:01:45.29" lane="4" heatid="14005">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:49.80" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="589" eventid="19" swimtime="00:00:43.72" lane="4" heatid="19003" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="186" birthdate="2008-01-01" gender="F" lastname="Zschegner" firstname="Lucy" license="0">
              <RESULTS>
                <RESULT resultid="590" eventid="10" swimtime="00:04:39.83" lane="4" heatid="10001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:04.31" />
                    <SPLIT distance="200" swimtime="00:02:16.55" />
                    <SPLIT distance="300" swimtime="00:03:30.82" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="591" eventid="13" swimtime="00:02:13.31" lane="5" heatid="13004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:01.58" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="592" eventid="18" swimtime="00:00:56.99" lane="5" heatid="18002" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="188" birthdate="2009-01-01" gender="F" lastname="Naupold" firstname="Celina" license="0">
              <RESULTS>
                <RESULT resultid="594" eventid="1" swimtime="00:00:22.10" lane="4" heatid="1002" />
                <RESULT resultid="595" eventid="8" swimtime="00:00:55.84" lane="1" heatid="8009" />
                <RESULT resultid="596" eventid="11" swimtime="00:00:25.55" lane="5" heatid="11010" />
                <RESULT resultid="597" eventid="18" status="DSQ" swimtime="00:00:00.00" lane="4" heatid="18002" comment="aufgegeben nach 5m" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="189" birthdate="2009-01-01" gender="M" lastname="Heydel" firstname="Linus" license="0">
              <RESULTS>
                <RESULT resultid="598" eventid="2" swimtime="00:00:21.78" lane="7" heatid="2002" />
                <RESULT resultid="599" eventid="9" swimtime="00:00:53.56" lane="8" heatid="9007" />
                <RESULT resultid="601" eventid="14" swimtime="00:02:03.65" lane="4" heatid="14004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:58.47" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="602" eventid="17" swimtime="00:04:33.25" lane="1" heatid="17003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:01.81" />
                    <SPLIT distance="200" swimtime="00:02:13.69" />
                    <SPLIT distance="300" swimtime="00:03:26.23" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="603" eventid="19" swimtime="00:00:56.89" lane="4" heatid="19002" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="191" birthdate="2010-01-01" gender="F" lastname="Dieke" firstname="Emelie" license="0">
              <RESULTS>
                <RESULT resultid="605" eventid="3" swimtime="00:00:33.50" lane="2" heatid="3001" />
                <RESULT resultid="606" eventid="8" swimtime="00:01:19.99" lane="5" heatid="8006" />
                <RESULT resultid="607" eventid="11" swimtime="00:00:31.32" lane="7" heatid="11007" />
                <RESULT resultid="608" eventid="13" swimtime="00:02:46.80" lane="8" heatid="13006">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:17.99" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="192" birthdate="2010-01-01" gender="M" lastname="Schröters" firstname="Paul" license="0">
              <RESULTS>
                <RESULT resultid="609" eventid="4" swimtime="00:00:38.47" lane="2" heatid="4002" />
                <RESULT resultid="610" eventid="9" swimtime="00:01:15.02" lane="8" heatid="9003" />
                <RESULT resultid="611" eventid="12" swimtime="00:00:32.69" lane="2" heatid="12001" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="195" birthdate="2011-01-01" gender="F" lastname="Volger" firstname="Eva" license="0">
              <RESULTS>
                <RESULT resultid="617" eventid="8" status="DSQ" swimtime="00:01:13.80" lane="1" heatid="8005" comment="falscher Start" />
                <RESULT resultid="618" eventid="11" swimtime="00:00:33.21" lane="8" heatid="11005" />
                <RESULT resultid="619" eventid="13" swimtime="00:02:46.24" lane="4" heatid="13003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:18.29" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="196" birthdate="2011-01-01" gender="M" lastname="Wyczisk" firstname="Johann" license="0">
              <RESULTS>
                <RESULT resultid="620" eventid="4" swimtime="00:00:32.50" lane="6" heatid="4002" />
                <RESULT resultid="621" eventid="9" swimtime="00:01:06.78" lane="4" heatid="9004" />
                <RESULT resultid="622" eventid="14" swimtime="00:02:26.32" lane="2" heatid="14003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:09.88" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="623" eventid="17" swimtime="00:05:13.50" lane="2" heatid="17002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:13.59" />
                    <SPLIT distance="200" swimtime="00:02:36.20" />
                    <SPLIT distance="300" swimtime="00:03:57.67" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="197" birthdate="2011-01-01" gender="F" lastname="Leonhardt" firstname="Ronja" license="0">
              <RESULTS>
                <RESULT resultid="624" eventid="8" swimtime="00:01:12.11" lane="6" heatid="8005" />
                <RESULT resultid="625" eventid="11" swimtime="00:00:33.52" lane="1" heatid="11005" />
                <RESULT resultid="626" eventid="13" swimtime="00:02:48.41" lane="2" heatid="13005">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:21.64" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="627" eventid="16" swimtime="00:05:50.95" lane="5" heatid="16002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:21.26" />
                    <SPLIT distance="200" swimtime="00:02:53.57" />
                    <SPLIT distance="300" swimtime="00:05:27.04" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="202" birthdate="2012-01-01" gender="M" lastname="Sochynskyi" firstname="Vadym" license="0">
              <RESULTS>
                <RESULT resultid="635" eventid="6" swimtime="00:00:33.39" lane="3" heatid="6002" />
                <RESULT resultid="636" eventid="9" swimtime="00:01:14.36" lane="7" heatid="9004" />
                <RESULT resultid="637" eventid="12" swimtime="00:00:33.38" lane="7" heatid="12003" />
                <RESULT resultid="638" eventid="14" swimtime="00:02:43.53" lane="3" heatid="14002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:18.63" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="639" eventid="17" swimtime="00:05:53.54" lane="1" heatid="17002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:20.26" />
                    <SPLIT distance="200" swimtime="00:02:52.88" />
                    <SPLIT distance="300" swimtime="00:04:24.59" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="203" birthdate="2013-01-01" gender="F" lastname="Jutzenka" firstname="Leonie" license="0">
              <RESULTS>
                <RESULT resultid="640" eventid="5" swimtime="00:00:44.34" lane="7" heatid="5002" />
                <RESULT resultid="641" eventid="8" swimtime="00:01:27.67" lane="7" heatid="8003" />
                <RESULT resultid="642" eventid="11" status="DSQ" swimtime="00:00:38.22" lane="5" heatid="11002" comment="falscher Start " />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="204" birthdate="2013-01-01" gender="M" lastname="Robenz" firstname="Ronny Jason" license="0">
              <RESULTS>
                <RESULT resultid="643" eventid="6" status="DSQ" swimtime="00:00:43.09" lane="2" heatid="6002" comment="falscher Stil bei 4m und 30m" />
                <RESULT resultid="644" eventid="9" swimtime="00:01:18.74" lane="5" heatid="9002" />
                <RESULT resultid="645" eventid="12" swimtime="00:00:33.76" lane="3" heatid="12002" />
                <RESULT resultid="646" eventid="14" swimtime="00:02:55.11" lane="8" heatid="14002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:24.63" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="205" birthdate="2014-01-01" gender="F" lastname="Zeil" firstname="Johanna" license="0">
              <RESULTS>
                <RESULT resultid="647" eventid="8" status="DSQ" swimtime="00:01:52.92" lane="8" heatid="8002" comment="falscher Start" />
                <RESULT resultid="648" eventid="11" swimtime="00:00:49.32" lane="4" heatid="11001" />
                <RESULT resultid="649" eventid="13" swimtime="00:04:12.58" lane="6" heatid="13002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:02:01.37" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="206" birthdate="2014-01-01" gender="F" lastname="Löffler" firstname="Leonie" license="0">
              <RESULTS>
                <RESULT resultid="650" eventid="8" swimtime="00:01:47.20" lane="4" heatid="8001" />
                <RESULT resultid="651" eventid="11" swimtime="00:00:42.90" lane="1" heatid="11002" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="207" birthdate="2014-01-01" gender="F" lastname="Blei" firstname="Lina" license="0">
              <RESULTS>
                <RESULT resultid="652" eventid="8" swimtime="00:01:46.50" lane="7" heatid="8002" />
                <RESULT resultid="653" eventid="11" swimtime="00:00:44.98" lane="7" heatid="11002" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="209" birthdate="2014-01-01" gender="M" lastname="Volger" firstname="Tom" license="0">
              <RESULTS>
                <RESULT resultid="655" eventid="6" swimtime="00:00:39.68" lane="7" heatid="6002" />
                <RESULT resultid="656" eventid="9" swimtime="00:01:20.42" lane="3" heatid="9003" />
                <RESULT resultid="657" eventid="12" swimtime="00:00:36.61" lane="6" heatid="12002" />
                <RESULT resultid="658" eventid="14" status="DSQ" swimtime="00:02:55.81" lane="6" heatid="14001" comment="falscher Start">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:25.57" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="210" birthdate="2015-01-01" gender="M" lastname="Viehhäuser" firstname="Aiden" license="0">
              <RESULTS>
                <RESULT resultid="659" eventid="6" status="DSQ" swimtime="00:00:53.32" lane="5" heatid="6001" comment="falscher Stil bei 2-10m" />
                <RESULT resultid="660" eventid="9" swimtime="00:01:36.12" lane="7" heatid="9002" />
                <RESULT resultid="661" eventid="12" swimtime="00:00:42.92" lane="6" heatid="12001" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="211" birthdate="2015-01-01" gender="F" lastname="Dieke" firstname="Anna" license="0">
              <RESULTS>
                <RESULT resultid="662" eventid="8" swimtime="00:01:40.51" lane="2" heatid="8002" />
                <RESULT resultid="663" eventid="11" swimtime="00:00:40.54" lane="2" heatid="11002" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="212" birthdate="2015-01-01" gender="M" lastname="Schulze" firstname="Joshua" license="0">
              <RESULTS>
                <RESULT resultid="664" eventid="6" swimtime="00:00:47.85" lane="3" heatid="6001" />
                <RESULT resultid="665" eventid="9" status="DSQ" swimtime="00:01:36.83" lane="3" heatid="9002" comment="falscher Start" />
                <RESULT resultid="666" eventid="12" swimtime="00:00:45.51" lane="4" heatid="12001" />
                <RESULT resultid="667" eventid="14" swimtime="00:03:29.01" lane="7" heatid="14001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:44.07" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="213" birthdate="2016-01-01" gender="F" lastname="Volger" firstname="Lea" license="0">
              <RESULTS>
                <RESULT resultid="668" eventid="5" status="DSQ" swimtime="00:00:46.55" lane="2" heatid="5002" comment="falscher Stil bei 40m" />
                <RESULT resultid="669" eventid="8" swimtime="00:01:33.72" lane="3" heatid="8002" />
                <RESULT resultid="670" eventid="11" swimtime="00:00:41.82" lane="6" heatid="11002" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="215" birthdate="2016-01-01" gender="M" lastname="Hierold" firstname="Theodor" license="0">
              <RESULTS>
                <RESULT resultid="672" eventid="6" swimtime="00:00:50.37" lane="4" heatid="6001" />
                <RESULT resultid="673" eventid="9" swimtime="00:01:33.52" lane="2" heatid="9002" />
                <RESULT resultid="674" eventid="12" swimtime="00:00:40.57" lane="1" heatid="12001" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY number="1" gender="M" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="593" eventid="21" swimtime="00:03:38.82" lane="8" heatid="21002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:53.96" />
                    <SPLIT distance="200" swimtime="00:01:55.03" />
                    <SPLIT distance="300" swimtime="00:02:54.18" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="189" number="1" />
                    <RELAYPOSITION athleteid="183" number="2" />
                    <RELAYPOSITION athleteid="184" number="3" />
                    <RELAYPOSITION athleteid="185" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" gender="F" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="604" eventid="20" status="WDR" swimtime="00:00:00.00" lane="7" heatid="20002">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="198" number="1" />
                    <RELAYPOSITION athleteid="197" number="2" />
                    <RELAYPOSITION athleteid="191" number="3" />
                    <RELAYPOSITION athleteid="188" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" gender="X" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="634" eventid="15" swimtime="00:02:29.04" lane="6" heatid="15001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:12.95" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="202" number="1" />
                    <RELAYPOSITION athleteid="203" number="2" />
                    <RELAYPOSITION athleteid="206" number="3" />
                    <RELAYPOSITION athleteid="204" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" gender="X" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="654" eventid="15" swimtime="00:03:00.40" lane="7" heatid="15001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:32.98" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="212" number="1" />
                    <RELAYPOSITION athleteid="207" number="2" />
                    <RELAYPOSITION athleteid="205" number="3" />
                    <RELAYPOSITION athleteid="209" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" gender="X" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="671" eventid="15" swimtime="00:02:56.71" lane="1" heatid="15001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:25.10" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="215" number="1" />
                    <RELAYPOSITION athleteid="213" number="2" />
                    <RELAYPOSITION athleteid="211" number="3" />
                    <RELAYPOSITION athleteid="210" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB name="TC fez Berlin" nation="GER" region="21" code="0">
          <ATHLETES>
            <ATHLETE athleteid="39" birthdate="2005-01-01" gender="F" lastname="Gawenda" firstname="Lara" license="0">
              <RESULTS>
                <RESULT resultid="171" eventid="1" swimtime="00:00:19.17" lane="6" heatid="1007" />
                <RESULT resultid="140" eventid="8" swimtime="00:00:45.28" lane="5" heatid="8014" />
                <RESULT resultid="180" eventid="11" swimtime="00:00:20.65" lane="5" heatid="11014" />
                <RESULT resultid="155" eventid="13" swimtime="00:01:42.89" lane="3" heatid="13011">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:50.13" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="163" eventid="16" swimtime="00:03:45.73" lane="4" heatid="16008">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:52.61" />
                    <SPLIT distance="200" swimtime="00:01:49.49" />
                    <SPLIT distance="300" swimtime="00:02:48.35" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="40" birthdate="2002-01-01" gender="F" lastname="Schikora" firstname="Johanna" license="0">
              <RESULTS>
                <RESULT resultid="172" eventid="1" swimtime="00:00:20.04" lane="4" heatid="1006" />
                <RESULT resultid="141" eventid="8" swimtime="00:00:45.99" lane="3" heatid="8014" />
                <RESULT resultid="168" eventid="10" swimtime="00:03:40.41" lane="2" heatid="10003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:53.65" />
                    <SPLIT distance="200" swimtime="00:01:49.97" />
                    <SPLIT distance="300" swimtime="00:02:45.72" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="154" eventid="13" swimtime="00:01:39.35" lane="5" heatid="13011">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:49.22" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="150" eventid="18" swimtime="00:00:47.03" lane="7" heatid="18005" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="41" birthdate="2007-01-01" gender="F" lastname="Schikora" firstname="Luise" license="0">
              <RESULTS>
                <RESULT resultid="173" eventid="1" swimtime="00:00:21.18" lane="8" heatid="1005" />
                <RESULT resultid="142" eventid="8" swimtime="00:00:49.77" lane="6" heatid="8012" />
                <RESULT resultid="181" eventid="11" swimtime="00:00:22.12" lane="1" heatid="11013" />
                <RESULT resultid="159" eventid="13" swimtime="00:01:56.03" lane="5" heatid="13008">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:52.72" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="42" birthdate="2014-01-01" gender="F" lastname="Rüdiger" firstname="Henrikje" license="0">
              <RESULTS>
                <RESULT resultid="176" eventid="5" swimtime="00:00:36.51" lane="6" heatid="5003" />
                <RESULT resultid="143" eventid="8" swimtime="00:01:21.40" lane="3" heatid="8003" />
                <RESULT resultid="182" eventid="11" swimtime="00:00:35.82" lane="8" heatid="11004" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="43" birthdate="2013-01-01" gender="F" lastname="Volkert" firstname="Sophia" license="0">
              <RESULTS>
                <RESULT resultid="177" eventid="5" swimtime="00:00:38.86" lane="8" heatid="5003" />
                <RESULT resultid="144" eventid="8" swimtime="00:01:29.49" lane="5" heatid="8003" />
                <RESULT resultid="183" eventid="11" swimtime="00:00:37.49" lane="6" heatid="11003" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="44" birthdate="2015-01-01" gender="F" lastname="Just" firstname="Elsa" license="0">
              <RESULTS>
                <RESULT resultid="178" eventid="5" status="DNS" swimtime="00:00:00.00" lane="3" heatid="5002" />
                <RESULT resultid="145" eventid="8" swimtime="00:01:38.65" lane="1" heatid="8002" />
                <RESULT resultid="184" eventid="11" swimtime="00:00:41.67" lane="4" heatid="11002" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="45" birthdate="1996-01-01" gender="M" lastname="Schustek" firstname="Fabian" license="0">
              <RESULTS>
                <RESULT resultid="175" eventid="2" swimtime="00:00:17.92" lane="4" heatid="2004" />
                <RESULT resultid="146" eventid="9" swimtime="00:00:43.49" lane="8" heatid="9010" />
                <RESULT resultid="185" eventid="12" swimtime="00:00:19.60" lane="1" heatid="12009" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="46" birthdate="2002-01-01" gender="M" lastname="Lebeau" firstname="Remy" license="0">
              <RESULTS>
                <RESULT resultid="147" eventid="9" swimtime="00:00:42.80" lane="4" heatid="9009" />
                <RESULT resultid="160" eventid="14" swimtime="00:01:37.42" lane="5" heatid="14006">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:47.99" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="151" eventid="19" swimtime="00:00:41.89" lane="7" heatid="19004" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="47" birthdate="2006-01-01" gender="M" lastname="Schlobohm" firstname="Enrico" license="0">
              <RESULTS>
                <RESULT resultid="174" eventid="2" swimtime="00:00:18.26" lane="7" heatid="2005" />
                <RESULT resultid="148" eventid="9" swimtime="00:00:44.75" lane="4" heatid="9008" />
                <RESULT resultid="186" eventid="12" swimtime="00:00:20.13" lane="7" heatid="12008" />
                <RESULT resultid="162" eventid="14" swimtime="00:01:54.15" lane="3" heatid="14005">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:53.90" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="48" birthdate="2014-01-01" gender="M" lastname="Bowe" firstname="Constantin" license="0">
              <RESULTS>
                <RESULT resultid="179" eventid="6" status="DSQ" swimtime="00:00:43.58" lane="6" heatid="6002" comment="falscher Start" />
                <RESULT resultid="149" eventid="9" status="DSQ" swimtime="00:01:26.64" lane="4" heatid="9002" comment="falscher Start" />
                <RESULT resultid="187" eventid="12" swimtime="00:00:39.59" lane="8" heatid="12002" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="49" birthdate="2005-01-01" gender="F" lastname="Tesch" firstname="Florentine" license="0">
              <RESULTS>
                <RESULT resultid="188" eventid="7" swimtime="00:08:17.36" lane="6" heatid="7004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:56.99" />
                    <SPLIT distance="200" swimtime="00:01:59.10" />
                    <SPLIT distance="300" swimtime="00:03:01.88" />
                    <SPLIT distance="400" swimtime="00:04:04.80" />
                    <SPLIT distance="500" swimtime="00:05:08.51" />
                    <SPLIT distance="600" swimtime="00:06:13.19" />
                    <SPLIT distance="700" swimtime="00:07:17.18" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="156" eventid="13" swimtime="00:01:53.26" lane="5" heatid="13010">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:52.87" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="164" eventid="16" swimtime="00:04:05.00" lane="7" heatid="16008">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:56.16" />
                    <SPLIT distance="200" swimtime="00:01:59.06" />
                    <SPLIT distance="300" swimtime="00:03:03.00" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="152" eventid="22" swimtime="00:15:44.96" lane="4" heatid="22002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:57.33" />
                    <SPLIT distance="200" swimtime="00:01:59.75" />
                    <SPLIT distance="300" swimtime="00:03:02.97" />
                    <SPLIT distance="400" swimtime="00:04:05.79" />
                    <SPLIT distance="500" swimtime="00:05:08.56" />
                    <SPLIT distance="600" swimtime="00:06:11.59" />
                    <SPLIT distance="700" swimtime="00:07:15.05" />
                    <SPLIT distance="800" swimtime="00:08:17.88" />
                    <SPLIT distance="900" swimtime="00:09:19.66" />
                    <SPLIT distance="1000" swimtime="00:10:22.00" />
                    <SPLIT distance="1100" swimtime="00:11:24.94" />
                    <SPLIT distance="1200" swimtime="00:12:29.13" />
                    <SPLIT distance="1300" swimtime="00:13:34.25" />
                    <SPLIT distance="1400" swimtime="00:14:40.33" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="50" birthdate="2006-01-01" gender="F" lastname="Ahnert" firstname="Paula" license="0">
              <RESULTS>
                <RESULT resultid="189" eventid="7" swimtime="00:08:03.03" lane="3" heatid="7004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:56.39" />
                    <SPLIT distance="200" swimtime="00:01:56.39" />
                    <SPLIT distance="300" swimtime="00:02:57.55" />
                    <SPLIT distance="400" swimtime="00:03:58.44" />
                    <SPLIT distance="500" swimtime="00:04:59.62" />
                    <SPLIT distance="600" swimtime="00:06:01.90" />
                    <SPLIT distance="700" swimtime="00:07:03.45" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="157" eventid="13" swimtime="00:01:44.01" lane="4" heatid="13010">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:50.63" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="165" eventid="16" swimtime="00:03:52.62" lane="1" heatid="16008">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:55.37" />
                    <SPLIT distance="200" swimtime="00:01:54.43" />
                    <SPLIT distance="300" swimtime="00:02:54.26" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="153" eventid="22" swimtime="00:15:35.27" lane="5" heatid="22002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:57.21" />
                    <SPLIT distance="200" swimtime="00:01:59.16" />
                    <SPLIT distance="300" swimtime="00:03:01.97" />
                    <SPLIT distance="400" swimtime="00:04:05.31" />
                    <SPLIT distance="500" swimtime="00:05:08.57" />
                    <SPLIT distance="600" swimtime="00:06:11.72" />
                    <SPLIT distance="700" swimtime="00:07:15.05" />
                    <SPLIT distance="800" swimtime="00:08:18.29" />
                    <SPLIT distance="900" swimtime="00:09:20.83" />
                    <SPLIT distance="1000" swimtime="00:10:24.24" />
                    <SPLIT distance="1100" swimtime="00:11:27.13" />
                    <SPLIT distance="1200" swimtime="00:12:30.25" />
                    <SPLIT distance="1300" swimtime="00:13:33.02" />
                    <SPLIT distance="1400" swimtime="00:14:34.65" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="51" birthdate="2006-01-01" gender="F" lastname="Zobel" firstname="Juliane" license="0">
              <RESULTS>
                <RESULT resultid="191" eventid="7" swimtime="00:08:50.48" lane="7" heatid="7003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:00.74" />
                    <SPLIT distance="200" swimtime="00:02:07.50" />
                    <SPLIT distance="300" swimtime="00:03:16.18" />
                    <SPLIT distance="400" swimtime="00:04:25.11" />
                    <SPLIT distance="500" swimtime="00:05:34.15" />
                    <SPLIT distance="600" swimtime="00:06:42.53" />
                    <SPLIT distance="700" swimtime="00:07:50.23" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="158" eventid="13" swimtime="00:01:55.01" lane="8" heatid="13009">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:54.72" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="166" eventid="16" swimtime="00:04:16.75" lane="5" heatid="16006">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:59.97" />
                    <SPLIT distance="200" swimtime="00:02:07.24" />
                    <SPLIT distance="300" swimtime="00:03:14.19" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="310" birthdate="2005-01-01" gender="M" lastname="Kwauka" firstname="Kevin" license="0" />
          </ATHLETES>
          <RELAYS>
            <RELAY number="1" gender="M" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="169" eventid="21" status="EXH" swimtime="00:02:57.28" lane="4" heatid="21002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:43.34" />
                    <SPLIT distance="200" swimtime="00:01:29.39" />
                    <SPLIT distance="300" swimtime="00:02:15.49" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="45" number="1" />
                    <RELAYPOSITION athleteid="310" number="2" />
                    <RELAYPOSITION athleteid="47" number="3" />
                    <RELAYPOSITION athleteid="46" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" gender="X" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="170" eventid="15" swimtime="00:02:36.64" lane="5" heatid="15001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:16.46" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="42" number="1" />
                    <RELAYPOSITION athleteid="48" number="2" />
                    <RELAYPOSITION athleteid="43" number="3" />
                    <RELAYPOSITION athleteid="44" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB name="TC Harz" nation="GER" region="27" code="0">
          <ATHLETES>
            <ATHLETE athleteid="133" birthdate="2008-01-01" gender="F" lastname="Weißemborn" firstname="Marnie" license="0">
              <RESULTS>
                <RESULT resultid="445" eventid="1" swimtime="00:00:20.58" lane="6" heatid="1005" />
                <RESULT resultid="414" eventid="8" swimtime="00:00:48.16" lane="4" heatid="8012" />
                <RESULT resultid="456" eventid="11" swimtime="00:00:22.12" lane="6" heatid="11013" />
                <RESULT resultid="425" eventid="13" swimtime="00:01:48.37" lane="2" heatid="13010">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:53.06" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="439" eventid="16" swimtime="00:04:08.54" lane="1" heatid="16006">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:00.37" />
                    <SPLIT distance="200" swimtime="00:02:05.92" />
                    <SPLIT distance="300" swimtime="00:03:08.56" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="134" birthdate="2007-01-01" gender="F" lastname="von Gynz Rekowski" firstname="Sophie" license="0">
              <RESULTS>
                <RESULT resultid="446" eventid="1" swimtime="00:00:22.06" lane="2" heatid="1005" />
                <RESULT resultid="415" eventid="8" swimtime="00:00:52.94" lane="4" heatid="8011" />
                <RESULT resultid="457" eventid="11" swimtime="00:00:23.58" lane="7" heatid="11012" />
                <RESULT resultid="427" eventid="13" swimtime="00:02:04.33" lane="3" heatid="13008">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:00.13" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="440" eventid="16" swimtime="00:04:33.19" lane="5" heatid="16005">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:03.34" />
                    <SPLIT distance="200" swimtime="00:02:13.27" />
                    <SPLIT distance="300" swimtime="00:03:25.41" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="135" birthdate="2011-01-01" gender="F" lastname="Chyla" firstname="Emma" license="0">
              <RESULTS>
                <RESULT resultid="416" eventid="8" swimtime="00:01:16.05" lane="4" heatid="8005" />
                <RESULT resultid="459" eventid="11" swimtime="00:00:32.71" lane="3" heatid="11004" />
                <RESULT resultid="429" eventid="13" swimtime="00:03:01.03" lane="3" heatid="13004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:22.28" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="136" birthdate="2012-01-01" gender="F" lastname="Krzizak" firstname="Lana" license="0">
              <RESULTS>
                <RESULT resultid="452" eventid="5" swimtime="00:00:36.59" lane="3" heatid="5003" />
                <RESULT resultid="417" eventid="8" swimtime="00:01:26.74" lane="8" heatid="8005" />
                <RESULT resultid="458" eventid="11" status="DSQ" swimtime="00:00:34.68" lane="6" heatid="11005" comment="falscher Start" />
                <RESULT resultid="432" eventid="13" swimtime="00:03:19.26" lane="1" heatid="13003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:35.46" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="137" birthdate="2012-01-01" gender="F" lastname="Dieck" firstname="Franziska" license="0">
              <RESULTS>
                <RESULT resultid="453" eventid="5" swimtime="00:00:35.50" lane="2" heatid="5003" />
                <RESULT resultid="418" eventid="8" swimtime="00:01:20.71" lane="1" heatid="8004" />
                <RESULT resultid="461" eventid="11" swimtime="00:00:33.81" lane="4" heatid="11003" />
                <RESULT resultid="431" eventid="13" swimtime="00:03:03.81" lane="5" heatid="13003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:27.48" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="138" birthdate="2011-01-01" gender="F" lastname="Dachner" firstname="Helena" license="0">
              <RESULTS>
                <RESULT resultid="419" eventid="8" swimtime="00:01:22.13" lane="8" heatid="8004" />
                <RESULT resultid="460" eventid="11" swimtime="00:00:34.36" lane="7" heatid="11004" />
                <RESULT resultid="430" eventid="13" swimtime="00:03:04.90" lane="2" heatid="13004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:30.46" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="139" birthdate="2008-01-01" gender="M" lastname="Härter" firstname="Fynn" license="0">
              <RESULTS>
                <RESULT resultid="451" eventid="2" swimtime="00:00:21.00" lane="2" heatid="2003" />
                <RESULT resultid="420" eventid="9" status="DSQ" swimtime="00:00:51.13" lane="2" heatid="9007" comment="falscher Start" />
                <RESULT resultid="464" eventid="12" swimtime="00:00:22.50" lane="6" heatid="12006" />
                <RESULT resultid="433" eventid="14" swimtime="00:01:54.85" lane="7" heatid="14005">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:54.78" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="441" eventid="17" swimtime="00:04:14.42" lane="2" heatid="17003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:56.53" />
                    <SPLIT distance="200" swimtime="00:02:04.37" />
                    <SPLIT distance="300" swimtime="00:03:12.76" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="140" birthdate="2013-01-01" gender="M" lastname="Hoffmeister" firstname="Oskar" license="0">
              <RESULTS>
                <RESULT resultid="454" eventid="6" swimtime="00:00:33.40" lane="4" heatid="6002" />
                <RESULT resultid="421" eventid="9" swimtime="00:01:10.65" lane="6" heatid="9004" />
                <RESULT resultid="467" eventid="12" swimtime="00:00:31.63" lane="1" heatid="12003" />
                <RESULT resultid="436" eventid="14" swimtime="00:02:34.80" lane="5" heatid="14001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:13.05" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="141" birthdate="2011-01-01" gender="M" lastname="Beier" firstname="Anton" license="0">
              <RESULTS>
                <RESULT resultid="422" eventid="9" swimtime="00:01:10.57" lane="8" heatid="9004" />
                <RESULT resultid="465" eventid="12" swimtime="00:00:30.29" lane="3" heatid="12003" />
                <RESULT resultid="435" eventid="14" status="DSQ" swimtime="00:02:33.40" lane="6" heatid="14002" comment="falsche Wende bei 150m ">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:12.84" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="142" birthdate="2009-01-01" gender="M" lastname="Piorun" firstname="Tariqe" license="0">
              <RESULTS>
                <RESULT resultid="423" eventid="9" status="DSQ" swimtime="00:01:05.92" lane="5" heatid="9003" comment="falscher Start" />
                <RESULT resultid="466" eventid="12" swimtime="00:00:30.18" lane="2" heatid="12003" />
                <RESULT resultid="434" eventid="14" swimtime="00:02:37.12" lane="5" heatid="14002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:16.02" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="143" birthdate="2012-01-01" gender="M" lastname="Neumann" firstname="Erik" license="0">
              <RESULTS>
                <RESULT resultid="455" eventid="6" swimtime="00:00:37.47" lane="5" heatid="6002" />
                <RESULT resultid="424" eventid="9" swimtime="00:01:11.06" lane="7" heatid="9003" />
                <RESULT resultid="468" eventid="12" swimtime="00:00:33.01" lane="2" heatid="12002" />
                <RESULT resultid="437" eventid="14" status="DSQ" swimtime="00:02:46.85" lane="3" heatid="14001" comment="Tauchzüge bei ca. 20-30m">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:26.25" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="144" birthdate="2007-01-01" gender="F" lastname="Risse" firstname="Elisabeth" license="0">
              <RESULTS>
                <RESULT resultid="447" eventid="1" swimtime="00:00:21.98" lane="1" heatid="1005" />
                <RESULT resultid="469" eventid="7" status="DSQ" swimtime="00:09:08.83" lane="2" heatid="7003" comment="15m nach Start übertaucht">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:56.99" />
                    <SPLIT distance="200" swimtime="00:02:03.98" />
                    <SPLIT distance="300" swimtime="00:03:13.01" />
                    <SPLIT distance="400" swimtime="00:04:24.05" />
                    <SPLIT distance="500" swimtime="00:05:35.97" />
                    <SPLIT distance="600" swimtime="00:06:48.69" />
                    <SPLIT distance="700" swimtime="00:08:00.53" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="426" eventid="13" swimtime="00:01:58.39" lane="3" heatid="13009">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:53.74" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="438" eventid="16" swimtime="00:04:24.23" lane="8" heatid="16007">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:57.86" />
                    <SPLIT distance="200" swimtime="00:02:05.08" />
                    <SPLIT distance="300" swimtime="00:03:15.43" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="145" birthdate="2009-01-01" gender="F" lastname="Zündel" firstname="Marlene" license="0">
              <RESULTS>
                <RESULT resultid="448" eventid="1" swimtime="00:00:24.38" lane="3" heatid="1003" />
                <RESULT resultid="470" eventid="7" swimtime="00:10:14.84" lane="3" heatid="7002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:05.53" />
                    <SPLIT distance="200" swimtime="00:02:22.24" />
                    <SPLIT distance="300" swimtime="00:02:40.18" />
                    <SPLIT distance="400" swimtime="00:05:00.27" />
                    <SPLIT distance="500" swimtime="00:06:19.65" />
                    <SPLIT distance="600" swimtime="00:07:41.83" />
                    <SPLIT distance="700" swimtime="00:08:59.49" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="428" eventid="13" swimtime="00:02:04.61" lane="6" heatid="13008">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:59.49" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="149" birthdate="2003-01-01" gender="M" lastname="Dalichow" firstname="Noah" license="0">
              <RESULTS>
                <RESULT resultid="449" eventid="2" swimtime="00:00:16.73" lane="2" heatid="2005" />
                <RESULT resultid="463" eventid="12" swimtime="00:00:19.73" lane="8" heatid="12008" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="150" birthdate="2004-01-01" gender="M" lastname="Hass" firstname="Jan Henrik" license="0">
              <RESULTS>
                <RESULT resultid="450" eventid="2" swimtime="00:00:18.25" lane="7" heatid="2004" />
                <RESULT resultid="462" eventid="12" swimtime="00:00:20.66" lane="1" heatid="12008" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY number="1" gender="F" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="442" eventid="20" swimtime="00:03:30.40" lane="6" heatid="20003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:51.49" />
                    <SPLIT distance="200" swimtime="00:01:46.10" />
                    <SPLIT distance="300" swimtime="00:02:36.85" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="133" number="1" />
                    <RELAYPOSITION athleteid="145" number="2" />
                    <RELAYPOSITION athleteid="144" number="3" />
                    <RELAYPOSITION athleteid="134" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" gender="F" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="443" eventid="20" swimtime="00:05:27.09" lane="5" heatid="20001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:17.68" />
                    <SPLIT distance="200" swimtime="00:02:38.17" />
                    <SPLIT distance="300" swimtime="00:04:01.67" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="135" number="1" />
                    <RELAYPOSITION athleteid="137" number="2" />
                    <RELAYPOSITION athleteid="138" number="3" />
                    <RELAYPOSITION athleteid="136" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" gender="M" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="444" eventid="21" swimtime="00:04:50.02" lane="1" heatid="21001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:12.48" />
                    <SPLIT distance="200" swimtime="00:02:22.09" />
                    <SPLIT distance="300" swimtime="00:03:38.78" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="141" number="1" />
                    <RELAYPOSITION athleteid="142" number="2" />
                    <RELAYPOSITION athleteid="143" number="3" />
                    <RELAYPOSITION athleteid="140" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB name="TC Marzahn e.V." nation="GER" region="21" code="0">
          <ATHLETES>
            <ATHLETE athleteid="266" birthdate="1965-01-01" gender="M" lastname="Ritzer" firstname="Andre" license="0">
              <RESULTS>
                <RESULT resultid="818" eventid="2" swimtime="00:00:23.47" lane="6" heatid="2002" />
                <RESULT resultid="819" eventid="9" swimtime="00:00:59.27" lane="5" heatid="9005" />
                <RESULT resultid="820" eventid="12" swimtime="00:00:26.36" lane="2" heatid="12005" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="267" birthdate="1971-01-01" gender="M" lastname="Tech" firstname="Matthias" license="0">
              <RESULTS>
                <RESULT resultid="821" eventid="2" swimtime="00:00:20.75" lane="1" heatid="2003" />
                <RESULT resultid="822" eventid="12" swimtime="00:00:23.60" lane="8" heatid="12006" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="269" birthdate="1977-01-01" gender="F" lastname="Lopez" firstname="Annett" license="0">
              <RESULTS>
                <RESULT resultid="824" eventid="8" swimtime="00:00:58.91" lane="3" heatid="8010" />
                <RESULT resultid="825" eventid="11" swimtime="00:00:26.10" lane="6" heatid="11010" />
                <RESULT resultid="826" eventid="13" swimtime="00:02:04.90" lane="4" heatid="13008">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:00.07" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="270" birthdate="1982-01-01" gender="F" lastname="Heilek" firstname="Sarah" license="0">
              <RESULTS>
                <RESULT resultid="827" eventid="8" swimtime="00:01:04.44" lane="4" heatid="8007" />
                <RESULT resultid="828" eventid="11" swimtime="00:00:29.37" lane="4" heatid="11007" />
                <RESULT resultid="829" eventid="13" swimtime="00:02:27.00" lane="7" heatid="13006">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:07.79" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="830" eventid="16" swimtime="00:05:39.49" lane="1" heatid="16004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:16.96" />
                    <SPLIT distance="200" swimtime="00:02:45.32" />
                    <SPLIT distance="300" swimtime="00:04:14.43" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="272" birthdate="2001-01-01" gender="M" lastname="Lopez" firstname="Marvin" license="0">
              <RESULTS>
                <RESULT resultid="832" eventid="2" swimtime="00:00:17.47" lane="6" heatid="2005" />
                <RESULT resultid="833" eventid="9" swimtime="00:00:43.54" lane="6" heatid="9009" />
                <RESULT resultid="834" eventid="12" swimtime="00:00:19.06" lane="7" heatid="12009" />
                <RESULT resultid="835" eventid="14" swimtime="00:01:42.05" lane="2" heatid="14006">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:49.00" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="274" birthdate="2005-01-01" gender="M" lastname="Kwauka" firstname="Kevin" license="0">
              <RESULTS>
                <RESULT resultid="840" eventid="2" swimtime="00:00:18.75" lane="3" heatid="2004" />
                <RESULT resultid="841" eventid="9" swimtime="00:00:45.38" lane="5" heatid="9008" />
                <RESULT resultid="842" eventid="12" swimtime="00:00:19.78" lane="2" heatid="12008" />
                <RESULT resultid="843" eventid="19" swimtime="00:00:44.68" lane="2" heatid="19003" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="276" birthdate="2005-01-01" gender="F" lastname="Eweleit" firstname="Laura" license="0">
              <RESULTS>
                <RESULT resultid="845" eventid="1" swimtime="00:00:18.96" lane="1" heatid="1007" />
                <RESULT resultid="955" eventid="7" swimtime="00:08:10.94" lane="7" heatid="7004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:56.02" />
                    <SPLIT distance="200" swimtime="00:01:57.12" />
                    <SPLIT distance="300" swimtime="00:02:59.90" />
                    <SPLIT distance="400" swimtime="00:04:02.87" />
                    <SPLIT distance="500" swimtime="00:05:06.50" />
                    <SPLIT distance="600" swimtime="00:06:09.99" />
                    <SPLIT distance="700" swimtime="00:07:11.58" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="846" eventid="8" swimtime="00:00:48.59" lane="6" heatid="8014" />
                <RESULT resultid="847" eventid="11" swimtime="00:00:21.08" lane="3" heatid="11014" />
                <RESULT resultid="848" eventid="16" swimtime="00:03:48.04" lane="3" heatid="16008">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:53.66" />
                    <SPLIT distance="200" swimtime="00:01:52.51" />
                    <SPLIT distance="300" swimtime="00:02:51.98" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="277" birthdate="2007-01-01" gender="F" lastname="Götz" firstname="Zoe" license="0">
              <RESULTS>
                <RESULT resultid="849" eventid="8" swimtime="00:00:52.57" lane="2" heatid="8012" />
                <RESULT resultid="850" eventid="11" swimtime="00:00:22.99" lane="8" heatid="11013" />
                <RESULT resultid="851" eventid="13" swimtime="00:02:00.15" lane="2" heatid="13009">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:58.06" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="852" eventid="18" swimtime="00:00:55.51" lane="2" heatid="18003" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="279" birthdate="2008-01-01" gender="F" lastname="Demmrich" firstname="Ella" license="0">
              <RESULTS>
                <RESULT resultid="854" eventid="1" swimtime="00:00:25.44" lane="1" heatid="1003" />
                <RESULT resultid="855" eventid="8" swimtime="00:01:01.07" lane="4" heatid="8009" />
                <RESULT resultid="856" eventid="11" swimtime="00:00:27.70" lane="3" heatid="11009" />
                <RESULT resultid="857" eventid="13" swimtime="00:02:13.41" lane="7" heatid="13007">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:02.89" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="858" eventid="16" swimtime="00:04:53.64" lane="1" heatid="16005">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:08.73" />
                    <SPLIT distance="200" swimtime="00:02:24.23" />
                    <SPLIT distance="300" swimtime="00:03:40.35" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="280" birthdate="2010-01-01" gender="F" lastname="Liedloff" firstname="Amelie" license="0">
              <RESULTS>
                <RESULT resultid="859" eventid="7" swimtime="00:10:39.41" lane="1" heatid="7003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:02.57" />
                    <SPLIT distance="200" swimtime="00:02:18.40" />
                    <SPLIT distance="300" swimtime="00:03:37.01" />
                    <SPLIT distance="400" swimtime="00:04:56.08" />
                    <SPLIT distance="500" swimtime="00:06:22.99" />
                    <SPLIT distance="600" swimtime="00:07:48.39" />
                    <SPLIT distance="700" swimtime="00:09:12.95" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="860" eventid="8" swimtime="00:00:54.46" lane="7" heatid="8012" />
                <RESULT resultid="861" eventid="11" swimtime="00:00:24.16" lane="2" heatid="11012" />
                <RESULT resultid="862" eventid="13" swimtime="00:02:06.26" lane="1" heatid="13009">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:59.33" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="863" eventid="16" swimtime="00:04:32.34" lane="4" heatid="16006">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:01.62" />
                    <SPLIT distance="200" swimtime="00:02:10.66" />
                    <SPLIT distance="300" swimtime="00:03:24.91" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="281" birthdate="2010-01-01" gender="F" lastname="Haupt" firstname="Lena" license="0">
              <RESULTS>
                <RESULT resultid="864" eventid="8" swimtime="00:00:55.45" lane="4" heatid="8010" />
                <RESULT resultid="865" eventid="11" swimtime="00:00:25.51" lane="3" heatid="11010" />
                <RESULT resultid="866" eventid="13" swimtime="00:02:11.06" lane="5" heatid="13007">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:03.31" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="867" eventid="16" swimtime="00:04:48.79" lane="6" heatid="16005">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:07.85" />
                    <SPLIT distance="200" swimtime="00:02:22.33" />
                    <SPLIT distance="300" swimtime="00:03:37.53" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="282" birthdate="2011-01-01" gender="F" lastname="Eweleit" firstname="Lenja" license="0">
              <RESULTS>
                <RESULT resultid="868" eventid="8" swimtime="00:00:59.54" lane="1" heatid="8010" />
                <RESULT resultid="869" eventid="11" swimtime="00:00:26.95" lane="5" heatid="11009" />
                <RESULT resultid="870" eventid="13" swimtime="00:02:13.68" lane="1" heatid="13007">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:06.18" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="871" eventid="16" swimtime="00:04:56.91" lane="7" heatid="16005">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:11.40" />
                    <SPLIT distance="200" swimtime="00:02:29.55" />
                    <SPLIT distance="300" swimtime="00:03:47.49" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY number="2" gender="X" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="817" eventid="15" swimtime="00:01:46.48" lane="5" heatid="15002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:56.70" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="266" number="1" />
                    <RELAYPOSITION athleteid="270" number="2" />
                    <RELAYPOSITION athleteid="267" number="3" />
                    <RELAYPOSITION athleteid="269" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="3" gender="F" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="853" eventid="20" swimtime="00:03:54.18" lane="1" heatid="20003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:55.47" />
                    <SPLIT distance="200" swimtime="00:01:55.59" />
                    <SPLIT distance="300" swimtime="00:02:56.12" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="280" number="1" />
                    <RELAYPOSITION athleteid="282" number="2" />
                    <RELAYPOSITION athleteid="279" number="3" />
                    <RELAYPOSITION athleteid="281" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB name="TC Potsdam e.V." nation="GER" region="19" code="0">
          <ATHLETES>
            <ATHLETE athleteid="85" birthdate="2003-01-01" gender="F" lastname="Junghans" firstname="Chiara" license="0">
              <RESULTS>
                <RESULT resultid="289" eventid="1" swimtime="00:00:19.88" lane="5" heatid="1005" />
                <RESULT resultid="279" eventid="8" swimtime="00:00:47.74" lane="3" heatid="8013" />
                <RESULT resultid="291" eventid="11" swimtime="00:00:21.66" lane="2" heatid="11013" />
                <RESULT resultid="286" eventid="16" swimtime="00:03:52.28" lane="6" heatid="16008">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:54.22" />
                    <SPLIT distance="200" swimtime="00:01:52.83" />
                    <SPLIT distance="300" swimtime="00:02:53.09" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="86" birthdate="1997-01-01" gender="F" lastname="Starke" firstname="Juliane" license="0">
              <RESULTS>
                <RESULT resultid="280" eventid="8" swimtime="00:00:47.34" lane="2" heatid="8013" />
                <RESULT resultid="283" eventid="13" swimtime="00:01:45.48" lane="6" heatid="13010">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:51.86" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="287" eventid="16" swimtime="00:03:47.41" lane="5" heatid="16007">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:54.00" />
                    <SPLIT distance="200" swimtime="00:01:52.60" />
                    <SPLIT distance="300" swimtime="00:02:51.90" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="87" birthdate="2011-01-01" gender="F" lastname="Oehme" firstname="Lilli" license="0">
              <RESULTS>
                <RESULT resultid="281" eventid="8" swimtime="00:01:19.23" lane="7" heatid="8004" />
                <RESULT resultid="292" eventid="11" swimtime="00:00:34.41" lane="4" heatid="11004" />
                <RESULT resultid="284" eventid="13" swimtime="00:02:59.23" lane="7" heatid="13004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:22.67" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="88" birthdate="2015-01-01" gender="F" lastname="Killat" firstname="Anna" license="0">
              <RESULTS>
                <RESULT resultid="290" eventid="5" swimtime="00:00:40.89" lane="6" heatid="5002" />
                <RESULT resultid="282" eventid="8" swimtime="00:01:25.42" lane="5" heatid="8002" />
                <RESULT resultid="293" eventid="11" swimtime="00:00:34.61" lane="3" heatid="11003" />
                <RESULT resultid="285" eventid="13" swimtime="00:03:04.48" lane="4" heatid="13002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:25.62" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY number="1" gender="F" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="288" eventid="20" swimtime="00:04:31.25" lane="3" heatid="20002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:50.06" />
                    <SPLIT distance="200" swimtime="00:02:18.21" />
                    <SPLIT distance="300" swimtime="00:03:44.96" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="86" number="1" />
                    <RELAYPOSITION athleteid="88" number="2" />
                    <RELAYPOSITION athleteid="87" number="3" />
                    <RELAYPOSITION athleteid="85" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB name="Tc submarin Pößneck" nation="GER" region="35" code="0">
          <ATHLETES>
            <ATHLETE athleteid="64" birthdate="2007-01-01" gender="F" lastname="Näther" firstname="Emilia" license="0">
              <RESULTS>
                <RESULT resultid="258" eventid="1" swimtime="00:00:19.56" lane="5" heatid="1006" />
                <RESULT resultid="216" eventid="8" swimtime="00:00:50.21" lane="8" heatid="8014" />
                <RESULT resultid="262" eventid="11" swimtime="00:00:21.53" lane="7" heatid="11014" />
                <RESULT resultid="238" eventid="13" swimtime="00:02:10.25" lane="7" heatid="13010">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:00.78" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="232" eventid="18" swimtime="00:00:48.65" lane="5" heatid="18003" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="65" birthdate="2010-01-01" gender="F" lastname="Matthes" firstname="Sophie" license="0">
              <RESULTS>
                <RESULT resultid="277" eventid="3" swimtime="00:00:26.78" lane="5" heatid="3001" />
                <RESULT resultid="217" eventid="8" swimtime="00:01:01.13" lane="7" heatid="8009" />
                <RESULT resultid="263" eventid="11" swimtime="00:00:27.37" lane="1" heatid="11009" />
                <RESULT resultid="239" eventid="13" swimtime="00:02:25.97" lane="1" heatid="13006">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:12.96" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="230" eventid="18" swimtime="00:01:10.87" lane="1" heatid="18001" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="66" birthdate="2012-01-01" gender="F" lastname="Kraus" firstname="Letizia Marie" license="0">
              <RESULTS>
                <RESULT resultid="260" eventid="5" swimtime="00:00:29.35" lane="4" heatid="5003" />
                <RESULT resultid="218" eventid="8" swimtime="00:01:03.77" lane="8" heatid="8007" />
                <RESULT resultid="264" eventid="11" swimtime="00:00:27.51" lane="3" heatid="11007" />
                <RESULT resultid="240" eventid="13" swimtime="00:02:21.17" lane="4" heatid="13005">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:07.13" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="249" eventid="16" swimtime="00:05:16.88" lane="2" heatid="16003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:08.95" />
                    <SPLIT distance="200" swimtime="00:02:33.57" />
                    <SPLIT distance="300" swimtime="00:03:59.47" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="67" birthdate="2011-01-01" gender="F" lastname="Müller" firstname="Emily" license="0">
              <RESULTS>
                <RESULT resultid="219" eventid="8" swimtime="00:01:08.26" lane="8" heatid="8006" />
                <RESULT resultid="265" eventid="11" swimtime="00:00:31.13" lane="8" heatid="11006" />
                <RESULT resultid="233" eventid="13" swimtime="00:02:37.93" lane="3" heatid="13001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:14.93" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="68" birthdate="2011-01-01" gender="F" lastname="Stenzel" firstname="Maja Lilou" license="0">
              <RESULTS>
                <RESULT resultid="220" eventid="8" swimtime="00:01:20.49" lane="4" heatid="8004" />
                <RESULT resultid="267" eventid="11" swimtime="00:00:34.71" lane="6" heatid="11004" />
                <RESULT resultid="235" eventid="13" swimtime="00:03:05.05" lane="2" heatid="13002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:32.09" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="69" birthdate="2013-01-01" gender="F" lastname="Huber" firstname="Sina" license="0">
              <RESULTS>
                <RESULT resultid="221" eventid="8" swimtime="00:01:14.30" lane="6" heatid="8004" />
                <RESULT resultid="266" eventid="11" swimtime="00:00:32.38" lane="3" heatid="11005" />
                <RESULT resultid="242" eventid="13" swimtime="00:02:52.10" lane="8" heatid="13003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:26.38" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="247" eventid="16" swimtime="00:06:17.09" lane="4" heatid="16001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:26.29" />
                    <SPLIT distance="200" swimtime="00:03:01.89" />
                    <SPLIT distance="300" swimtime="00:04:44.58" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="70" birthdate="2013-01-01" gender="F" lastname="Werner" firstname="Zoe" license="0">
              <RESULTS>
                <RESULT resultid="222" eventid="8" status="DNS" swimtime="00:00:00.00" lane="2" heatid="8004" />
                <RESULT resultid="270" eventid="11" swimtime="00:00:37.17" lane="2" heatid="11003" />
                <RESULT resultid="236" eventid="13" swimtime="00:03:05.75" lane="1" heatid="13002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:32.78" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="71" birthdate="2013-01-01" gender="F" lastname="Dietzel" firstname="Hanna" license="0">
              <RESULTS>
                <RESULT resultid="259" eventid="5" swimtime="00:00:46.60" lane="5" heatid="5001" />
                <RESULT resultid="223" eventid="8" swimtime="00:01:27.93" lane="2" heatid="8003" />
                <RESULT resultid="271" eventid="11" swimtime="00:00:36.65" lane="1" heatid="11003" />
                <RESULT resultid="234" eventid="13" status="DSQ" swimtime="00:03:18.66" lane="4" heatid="13001" comment="falscher Start">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:34.36" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="72" birthdate="2013-01-01" gender="F" lastname="Schmidt" firstname="Ylva" license="0">
              <RESULTS>
                <RESULT resultid="261" eventid="5" swimtime="00:00:40.29" lane="5" heatid="5003" />
                <RESULT resultid="224" eventid="8" swimtime="00:01:20.10" lane="1" heatid="8003" />
                <RESULT resultid="269" eventid="11" swimtime="00:00:36.42" lane="5" heatid="11003" />
                <RESULT resultid="241" eventid="13" swimtime="00:02:59.54" lane="7" heatid="13003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:24.36" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="73" birthdate="2013-01-01" gender="F" lastname="Trunk" firstname="Mila" license="0">
              <RESULTS>
                <RESULT resultid="225" eventid="8" swimtime="00:01:17.78" lane="6" heatid="8002" />
                <RESULT resultid="268" eventid="11" swimtime="00:00:35.60" lane="2" heatid="11004" />
                <RESULT resultid="246" eventid="16" swimtime="00:06:31.38" lane="1" heatid="16002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:31.48" />
                    <SPLIT distance="200" swimtime="00:03:15.09" />
                    <SPLIT distance="300" swimtime="00:04:56.36" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="74" birthdate="2013-01-01" gender="M" lastname="Langlotz" firstname="Lennert" license="0">
              <RESULTS>
                <RESULT resultid="226" eventid="9" swimtime="00:01:25.78" lane="4" heatid="9001" />
                <RESULT resultid="276" eventid="12" status="DSQ" swimtime="00:00:37.02" lane="3" heatid="12001" comment="fakscher Start" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="75" birthdate="2011-01-01" gender="M" lastname="Knoblich" firstname="Paul" license="0">
              <RESULTS>
                <RESULT resultid="278" eventid="4" swimtime="00:00:33.74" lane="5" heatid="4001" />
                <RESULT resultid="227" eventid="9" swimtime="00:01:14.57" lane="4" heatid="9003" />
                <RESULT resultid="273" eventid="12" swimtime="00:00:31.46" lane="4" heatid="12002" />
                <RESULT resultid="244" eventid="14" swimtime="00:02:46.40" lane="2" heatid="14002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:21.46" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="250" eventid="17" swimtime="00:06:03.18" lane="5" heatid="17001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:24.65" />
                    <SPLIT distance="200" swimtime="00:02:59.50" />
                    <SPLIT distance="300" swimtime="00:04:34.20" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="76" birthdate="2011-01-01" gender="M" lastname="Rattke" firstname="Carlos" license="0">
              <RESULTS>
                <RESULT resultid="228" eventid="9" swimtime="00:01:10.86" lane="6" heatid="9003" />
                <RESULT resultid="274" eventid="12" swimtime="00:00:32.84" lane="5" heatid="12002" />
                <RESULT resultid="245" eventid="14" swimtime="00:02:41.08" lane="7" heatid="14002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:22.08" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="77" birthdate="2013-01-01" gender="M" lastname="Dommler" firstname="Fabrice" license="0">
              <RESULTS>
                <RESULT resultid="229" eventid="9" swimtime="00:01:18.58" lane="1" heatid="9003" />
                <RESULT resultid="275" eventid="12" swimtime="00:00:34.38" lane="1" heatid="12002" />
                <RESULT resultid="243" eventid="14" swimtime="00:03:08.42" lane="1" heatid="14001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:33.98" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="78" birthdate="2005-01-01" gender="F" lastname="Heinze" firstname="Charlotte" license="0">
              <RESULTS>
                <RESULT resultid="257" eventid="1" swimtime="00:00:19.03" lane="8" heatid="1007" />
                <RESULT resultid="251" eventid="10" swimtime="00:04:01.19" lane="7" heatid="10002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:54.45" />
                    <SPLIT distance="200" swimtime="00:01:55.75" />
                    <SPLIT distance="300" swimtime="00:02:59.90" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="237" eventid="13" swimtime="00:01:54.18" lane="3" heatid="13010">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:54.22" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="231" eventid="18" swimtime="00:00:44.12" lane="4" heatid="18004" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="84" birthdate="2015-01-01" gender="F" lastname="Huber" firstname="Karla" license="0">
              <RESULTS>
                <RESULT resultid="272" eventid="11" swimtime="00:00:46.95" lane="8" heatid="11002" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY number="1" gender="F" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="252" eventid="20" swimtime="00:05:19.04" lane="6" heatid="20002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:21.43" />
                    <SPLIT distance="200" swimtime="00:02:44.42" />
                    <SPLIT distance="300" swimtime="00:04:10.46" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="69" number="1" />
                    <RELAYPOSITION athleteid="70" number="2" />
                    <RELAYPOSITION athleteid="73" number="3" />
                    <RELAYPOSITION athleteid="66" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" gender="F" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="253" eventid="20" swimtime="00:05:31.61" lane="3" heatid="20001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:25.18" />
                    <SPLIT distance="200" swimtime="00:02:58.18" />
                    <SPLIT distance="300" swimtime="00:04:20.47" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="68" number="1" />
                    <RELAYPOSITION athleteid="71" number="2" />
                    <RELAYPOSITION athleteid="72" number="3" />
                    <RELAYPOSITION athleteid="67" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" gender="M" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="254" eventid="21" swimtime="00:05:24.42" lane="8" heatid="21001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:12.24" />
                    <SPLIT distance="200" swimtime="00:02:42.47" />
                    <SPLIT distance="300" swimtime="00:04:09.16" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="76" number="1" />
                    <RELAYPOSITION athleteid="74" number="2" />
                    <RELAYPOSITION athleteid="77" number="3" />
                    <RELAYPOSITION athleteid="75" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" gender="X" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="255" eventid="15" swimtime="00:02:15.52" lane="4" heatid="15001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:10.82" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="69" number="1" />
                    <RELAYPOSITION athleteid="70" number="2" />
                    <RELAYPOSITION athleteid="73" number="3" />
                    <RELAYPOSITION athleteid="66" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" gender="X" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="256" eventid="15" swimtime="00:02:27.67" lane="2" heatid="15001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:13.15" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="71" number="1" />
                    <RELAYPOSITION athleteid="77" number="2" />
                    <RELAYPOSITION athleteid="74" number="3" />
                    <RELAYPOSITION athleteid="72" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB name="TSC Schwandorf e.V." nation="GER" region="34" code="0">
          <ATHLETES>
            <ATHLETE athleteid="31" birthdate="2010-01-01" gender="F" lastname="Seitz" firstname="Melina" license="0">
              <RESULTS>
                <RESULT resultid="121" eventid="8" swimtime="00:01:00.90" lane="6" heatid="8009" />
                <RESULT resultid="130" eventid="11" swimtime="00:00:27.45" lane="2" heatid="11009" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="32" birthdate="2011-01-01" gender="F" lastname="Maget" firstname="Matilda" license="0">
              <RESULTS>
                <RESULT resultid="122" eventid="8" status="DSQ" swimtime="00:01:06.67" lane="7" heatid="8007" comment="falscher Start" />
                <RESULT resultid="131" eventid="11" swimtime="00:00:29.23" lane="1" heatid="11008" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="33" birthdate="2007-01-01" gender="F" lastname="Böhner" firstname="Madeleine" license="0">
              <RESULTS>
                <RESULT resultid="123" eventid="8" swimtime="00:01:11.42" lane="2" heatid="8006" />
                <RESULT resultid="132" eventid="11" swimtime="00:00:31.74" lane="1" heatid="11006" />
                <RESULT resultid="125" eventid="18" swimtime="00:01:16.89" lane="6" heatid="18001" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="34" birthdate="2004-01-01" gender="F" lastname="Kohler" firstname="Nina" license="0">
              <RESULTS>
                <RESULT resultid="128" eventid="1" swimtime="00:00:18.18" lane="5" heatid="1007" />
                <RESULT resultid="129" eventid="11" swimtime="00:00:20.10" lane="4" heatid="11014" />
                <RESULT resultid="124" eventid="18" swimtime="00:00:41.94" lane="6" heatid="18005" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="35" birthdate="2007-01-01" gender="F" lastname="Rödl" firstname="Emily" license="0">
              <RESULTS>
                <RESULT resultid="133" eventid="7" swimtime="00:08:24.20" lane="4" heatid="7002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:56.38" />
                    <SPLIT distance="200" swimtime="00:01:59.61" />
                    <SPLIT distance="300" swimtime="00:03:05.12" />
                    <SPLIT distance="400" swimtime="00:04:10.47" />
                    <SPLIT distance="500" swimtime="00:05:15.36" />
                    <SPLIT distance="600" swimtime="00:06:20.63" />
                    <SPLIT distance="700" swimtime="00:07:24.29" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="126" eventid="16" swimtime="00:04:00.87" lane="2" heatid="16007">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:55.73" />
                    <SPLIT distance="200" swimtime="00:01:58.29" />
                    <SPLIT distance="300" swimtime="00:03:01.78" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY number="1" gender="F" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="127" eventid="20" swimtime="00:03:37.89" lane="7" heatid="20003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:44.51" />
                    <SPLIT distance="200" swimtime="00:01:49.75" />
                    <SPLIT distance="300" swimtime="00:02:50.51" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="34" number="1" />
                    <RELAYPOSITION athleteid="32" number="2" />
                    <RELAYPOSITION athleteid="31" number="3" />
                    <RELAYPOSITION athleteid="35" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB name="TSC Weimar e.V." nation="GER" region="35" code="0">
          <ATHLETES>
            <ATHLETE athleteid="90" birthdate="2012-01-01" gender="F" lastname="Riemann" firstname="Ada" license="0">
              <RESULTS>
                <RESULT resultid="348" eventid="5" swimtime="00:00:41.47" lane="8" heatid="5002" />
                <RESULT resultid="294" eventid="8" swimtime="00:01:26.65" lane="2" heatid="8001" />
                <RESULT resultid="355" eventid="11" swimtime="00:00:37.15" lane="5" heatid="11001" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="91" birthdate="2012-01-01" gender="F" lastname="Gollhardt" firstname="Fridoline" license="0">
              <RESULTS>
                <RESULT resultid="349" eventid="5" swimtime="00:00:39.13" lane="3" heatid="5001" />
                <RESULT resultid="295" eventid="8" swimtime="00:01:37.67" lane="6" heatid="8001" />
                <RESULT resultid="356" eventid="11" swimtime="00:00:34.42" lane="2" heatid="11001" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="92" birthdate="2013-01-01" gender="F" lastname="Erfurt" firstname="Marit" license="0">
              <RESULTS>
                <RESULT resultid="350" eventid="5" status="DSQ" swimtime="00:00:43.11" lane="1" heatid="5002" comment="falscher Stil bei 30m" />
                <RESULT resultid="296" eventid="8" swimtime="00:01:26.88" lane="3" heatid="8001" />
                <RESULT resultid="357" eventid="11" swimtime="00:00:40.08" lane="3" heatid="11001" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="94" birthdate="2010-01-01" gender="F" lastname="Pontes" firstname="Lena" license="0">
              <RESULTS>
                <RESULT resultid="298" eventid="8" swimtime="00:01:04.21" lane="3" heatid="8006" />
                <RESULT resultid="359" eventid="11" swimtime="00:00:26.92" lane="8" heatid="11007" />
                <RESULT resultid="321" eventid="13" swimtime="00:02:35.88" lane="8" heatid="13005">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:17.53" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="95" birthdate="2011-01-01" gender="F" lastname="Hüttig" firstname="Maline" license="0">
              <RESULTS>
                <RESULT resultid="299" eventid="8" swimtime="00:01:09.62" lane="2" heatid="8005" />
                <RESULT resultid="360" eventid="11" swimtime="00:00:28.30" lane="6" heatid="11006" />
                <RESULT resultid="322" eventid="13" swimtime="00:02:51.44" lane="1" heatid="13005">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:21.71" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="96" birthdate="2010-01-01" gender="F" lastname="Seyfarth" firstname="Anni" license="0">
              <RESULTS>
                <RESULT resultid="300" eventid="8" swimtime="00:01:04.83" lane="5" heatid="8004" />
                <RESULT resultid="361" eventid="11" swimtime="00:00:28.63" lane="4" heatid="11005" />
                <RESULT resultid="323" eventid="13" swimtime="00:02:27.18" lane="1" heatid="13004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:11.28" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="329" eventid="16" swimtime="00:05:30.99" lane="5" heatid="16001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:15.31" />
                    <SPLIT distance="200" swimtime="00:02:42.80" />
                    <SPLIT distance="300" swimtime="00:04:10.77" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="97" birthdate="2012-01-01" gender="F" lastname="Linne" firstname="Nora" license="0">
              <RESULTS>
                <RESULT resultid="351" eventid="5" swimtime="00:00:36.71" lane="4" heatid="5001" />
                <RESULT resultid="301" eventid="8" status="DSQ" swimtime="00:01:26.10" lane="6" heatid="8003" comment="falscher Start" />
                <RESULT resultid="362" eventid="11" swimtime="00:00:39.63" lane="8" heatid="11003" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="98" birthdate="2014-01-01" gender="M" lastname="Schmeißer" firstname="Edwin" license="0">
              <RESULTS>
                <RESULT resultid="354" eventid="6" status="DSQ" swimtime="00:00:43.54" lane="1" heatid="6002" comment="falscher Start" />
                <RESULT resultid="302" eventid="9" swimtime="00:01:33.15" lane="5" heatid="9001" />
                <RESULT resultid="375" eventid="12" status="DSQ" swimtime="00:00:45.09" lane="7" heatid="12001" comment="falscher Start" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="100" birthdate="2013-01-01" gender="M" lastname="Kröckel" firstname="Maximilian" license="0">
              <RESULTS>
                <RESULT resultid="304" eventid="9" status="DSQ" swimtime="00:01:38.83" lane="3" heatid="9001" comment="falscher Start" />
                <RESULT resultid="364" eventid="12" swimtime="00:00:46.41" lane="8" heatid="12001" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="101" birthdate="2005-01-01" gender="M" lastname="Linne" firstname="Georg" license="0">
              <RESULTS>
                <RESULT resultid="339" eventid="2" swimtime="00:00:17.50" lane="3" heatid="2005" />
                <RESULT resultid="305" eventid="9" swimtime="00:00:43.04" lane="8" heatid="9009" />
                <RESULT resultid="331" eventid="10" swimtime="00:03:16.53" lane="3" heatid="10003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:44.48" />
                    <SPLIT distance="200" swimtime="00:01:33.60" />
                    <SPLIT distance="300" swimtime="00:02:25.63" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="324" eventid="14" swimtime="00:01:38.09" lane="7" heatid="14006">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:47.40" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="315" eventid="19" swimtime="00:00:39.16" lane="2" heatid="19004" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="102" birthdate="2006-01-01" gender="M" lastname="Hauser" firstname="Theo" license="0">
              <RESULTS>
                <RESULT resultid="341" eventid="2" swimtime="00:00:19.22" lane="6" heatid="2004" />
                <RESULT resultid="306" eventid="9" swimtime="00:00:46.45" lane="6" heatid="9008" />
                <RESULT resultid="366" eventid="12" swimtime="00:00:19.89" lane="5" heatid="12007" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="103" birthdate="2004-01-01" gender="M" lastname="Röthlich" firstname="Nils" license="0">
              <RESULTS>
                <RESULT resultid="342" eventid="2" swimtime="00:00:19.55" lane="2" heatid="2004" />
                <RESULT resultid="307" eventid="9" swimtime="00:00:46.72" lane="7" heatid="9008" />
                <RESULT resultid="365" eventid="12" swimtime="00:00:21.00" lane="4" heatid="12007" />
                <RESULT resultid="316" eventid="19" swimtime="00:00:46.34" lane="6" heatid="19003" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="104" birthdate="2008-01-01" gender="M" lastname="Kraft" firstname="Simon" license="0">
              <RESULTS>
                <RESULT resultid="340" eventid="2" swimtime="00:00:18.18" lane="8" heatid="2005" />
                <RESULT resultid="308" eventid="9" swimtime="00:00:47.14" lane="4" heatid="9007" />
                <RESULT resultid="367" eventid="12" swimtime="00:00:20.55" lane="2" heatid="12007" />
                <RESULT resultid="317" eventid="19" swimtime="00:00:41.39" lane="7" heatid="19003" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="106" birthdate="2011-01-01" gender="M" lastname="Bellmann" firstname="Lennart" license="0">
              <RESULTS>
                <RESULT resultid="377" eventid="4" swimtime="00:00:27.76" lane="1" heatid="4002" />
                <RESULT resultid="310" eventid="9" swimtime="00:00:58.98" lane="8" heatid="9006" />
                <RESULT resultid="369" eventid="12" swimtime="00:00:25.70" lane="3" heatid="12005" />
                <RESULT resultid="325" eventid="14" swimtime="00:02:38.43" lane="7" heatid="14004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:15.02" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="320" eventid="19" swimtime="00:01:11.35" lane="8" heatid="19002" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="107" birthdate="2010-01-01" gender="M" lastname="Bellmann" firstname="Arvid" license="0">
              <RESULTS>
                <RESULT resultid="378" eventid="4" swimtime="00:00:26.35" lane="3" heatid="4002" />
                <RESULT resultid="311" eventid="9" swimtime="00:00:59.23" lane="7" heatid="9005" />
                <RESULT resultid="370" eventid="12" swimtime="00:00:26.13" lane="7" heatid="12005" />
                <RESULT resultid="327" eventid="14" swimtime="00:02:12.85" lane="4" heatid="14003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:04.71" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="319" eventid="19" swimtime="00:01:01.97" lane="1" heatid="19002" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="108" birthdate="2009-01-01" gender="M" lastname="Klabunde" firstname="Kalle" license="0">
              <RESULTS>
                <RESULT resultid="312" eventid="9" swimtime="00:01:03.33" lane="8" heatid="9005" />
                <RESULT resultid="373" eventid="12" swimtime="00:00:27.59" lane="8" heatid="12004" />
                <RESULT resultid="326" eventid="14" swimtime="00:02:22.58" lane="1" heatid="14004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:07.86" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="109" birthdate="1956-01-01" gender="M" lastname="Scheffzük" firstname="Olaf" license="0">
              <RESULTS>
                <RESULT resultid="345" eventid="2" swimtime="00:00:28.58" lane="5" heatid="2001" />
                <RESULT resultid="313" eventid="9" swimtime="00:01:00.69" lane="5" heatid="9004" />
                <RESULT resultid="372" eventid="12" swimtime="00:00:27.33" lane="4" heatid="12004" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="110" birthdate="2002-01-01" gender="F" lastname="Kluge" firstname="Paula" license="0">
              <RESULTS>
                <RESULT resultid="338" eventid="1" swimtime="00:00:18.84" lane="7" heatid="1007" />
                <RESULT resultid="332" eventid="10" swimtime="00:04:08.77" lane="7" heatid="10003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:49.65" />
                    <SPLIT distance="200" swimtime="00:01:54.16" />
                    <SPLIT distance="300" swimtime="00:03:02.52" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="358" eventid="11" swimtime="00:00:21.40" lane="1" heatid="11014" />
                <RESULT resultid="314" eventid="18" swimtime="00:00:43.32" lane="5" heatid="18005" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="111" birthdate="2002-01-01" gender="F" lastname="Stein" firstname="Franziska" license="0">
              <RESULTS>
                <RESULT resultid="330" eventid="16" swimtime="00:04:03.59" lane="8" heatid="16006">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:55.73" />
                    <SPLIT distance="200" swimtime="00:01:58.86" />
                    <SPLIT distance="300" swimtime="00:03:02.29" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="117" birthdate="1965-01-01" gender="M" lastname="Krieg" firstname="Marcus" license="0">
              <RESULTS>
                <RESULT resultid="344" eventid="2" swimtime="00:00:26.23" lane="8" heatid="2002" />
                <RESULT resultid="371" eventid="12" swimtime="00:00:26.00" lane="1" heatid="12005" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="118" birthdate="1960-01-01" gender="M" lastname="Kaleta" firstname="Bernd" license="0">
              <RESULTS>
                <RESULT resultid="346" eventid="2" swimtime="00:00:34.11" lane="6" heatid="2001" />
                <RESULT resultid="374" eventid="12" swimtime="00:00:31.02" lane="4" heatid="12003" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="119" birthdate="1973-01-01" gender="M" lastname="Brych" firstname="Ronald" license="0">
              <RESULTS>
                <RESULT resultid="347" eventid="2" swimtime="00:00:30.77" lane="2" heatid="2001" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="175" birthdate="1971-01-01" gender="F" lastname="Klabunde" firstname="Monique" license="0" />
            <ATHLETE athleteid="176" birthdate="1968-01-01" gender="M" lastname="Klabunde" firstname="Sven" license="0" />
            <ATHLETE athleteid="305" birthdate="1965-01-01" gender="M" lastname="Naue" firstname="Lutz" license="0" />
            <ATHLETE athleteid="306" birthdate="1967-01-01" gender="M" lastname="Wurzbacher" firstname="Markus" license="0" />
            <ATHLETE athleteid="309" birthdate="2004-01-01" gender="M" lastname="Haufe" firstname="Elias" license="0" />
          </ATHLETES>
          <RELAYS>
            <RELAY number="1" gender="M" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="333" eventid="21" swimtime="00:03:01.89" lane="2" heatid="21002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:43.72" />
                    <SPLIT distance="200" swimtime="00:01:30.48" />
                    <SPLIT distance="300" swimtime="00:02:16.08" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="101" number="1" />
                    <RELAYPOSITION athleteid="103" number="2" />
                    <RELAYPOSITION athleteid="104" number="3" />
                    <RELAYPOSITION athleteid="309" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" gender="X" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="334" eventid="21" swimtime="00:03:51.50" lane="5" heatid="21001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:54.85" />
                    <SPLIT distance="200" swimtime="00:01:55.43" />
                    <SPLIT distance="300" swimtime="00:02:54.55" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="175" number="1" />
                    <RELAYPOSITION athleteid="109" number="2" />
                    <RELAYPOSITION athleteid="117" number="3" />
                    <RELAYPOSITION athleteid="176" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" gender="M" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="335" eventid="21" status="DSQ" swimtime="00:04:23.57" lane="6" heatid="21001" comment="falscher Start">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:04.74" />
                    <SPLIT distance="200" swimtime="00:02:15.66" />
                    <SPLIT distance="300" swimtime="00:03:17.46" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="305" number="1" />
                    <RELAYPOSITION athleteid="118" number="2" />
                    <RELAYPOSITION athleteid="306" number="3" />
                    <RELAYPOSITION athleteid="119" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" gender="X" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="336" eventid="15" swimtime="00:02:33.49" lane="8" heatid="15001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:18.49" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="92" number="1" />
                    <RELAYPOSITION athleteid="90" number="2" />
                    <RELAYPOSITION athleteid="91" number="3" />
                    <RELAYPOSITION athleteid="97" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" gender="X" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="337" eventid="15" swimtime="00:01:42.69" lane="6" heatid="15002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:51.48" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="175" number="1" />
                    <RELAYPOSITION athleteid="109" number="2" />
                    <RELAYPOSITION athleteid="117" number="3" />
                    <RELAYPOSITION athleteid="176" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB name="TSG TU Ilmenau 56 e.V." nation="GER" region="35" code="0">
          <ATHLETES>
            <ATHLETE athleteid="285" birthdate="1998-01-01" gender="M" lastname="Rose" firstname="Jonas" license="0">
              <RESULTS>
                <RESULT resultid="875" eventid="7" swimtime="00:08:45.35" lane="5" heatid="7003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:57.99" />
                    <SPLIT distance="200" swimtime="00:02:03.21" />
                    <SPLIT distance="300" swimtime="00:03:09.96" />
                    <SPLIT distance="400" swimtime="00:04:17.23" />
                    <SPLIT distance="500" swimtime="00:05:24.82" />
                    <SPLIT distance="600" swimtime="00:06:33.89" />
                    <SPLIT distance="700" swimtime="00:07:42.60" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="876" eventid="10" swimtime="00:03:48.28" lane="1" heatid="10003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:50.12" />
                    <SPLIT distance="200" swimtime="00:01:48.46" />
                    <SPLIT distance="300" swimtime="00:02:47.51" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="877" eventid="19" swimtime="00:00:43.21" lane="5" heatid="19003" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="286" birthdate="2001-01-01" gender="M" lastname="Pohl" firstname="Enrico" license="0">
              <RESULTS>
                <RESULT resultid="878" eventid="2" swimtime="00:00:15.98" lane="3" heatid="2006" />
                <RESULT resultid="879" eventid="9" swimtime="00:00:40.02" lane="7" heatid="9010" />
                <RESULT resultid="880" eventid="12" swimtime="00:00:17.74" lane="6" heatid="12009" />
                <RESULT resultid="881" eventid="14" swimtime="00:01:45.01" lane="8" heatid="14006">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:48.78" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="287" birthdate="2004-01-01" gender="M" lastname="Dombrowsky" firstname="Lennard" license="0">
              <RESULTS>
                <RESULT resultid="883" eventid="7" swimtime="00:08:34.34" lane="8" heatid="7004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:53.16" />
                    <SPLIT distance="200" swimtime="00:01:58.40" />
                    <SPLIT distance="300" swimtime="00:03:02.62" />
                    <SPLIT distance="400" swimtime="00:04:08.39" />
                    <SPLIT distance="500" swimtime="00:05:15.18" />
                    <SPLIT distance="600" swimtime="00:06:22.81" />
                    <SPLIT distance="700" swimtime="00:07:28.30" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="884" eventid="9" swimtime="00:00:44.45" lane="1" heatid="9009" />
                <RESULT resultid="885" eventid="12" swimtime="00:00:20.02" lane="6" heatid="12008" />
                <RESULT resultid="886" eventid="14" swimtime="00:01:49.24" lane="1" heatid="14006">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:51.11" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="887" eventid="22" status="DSQ" swimtime="00:00:00.00" lane="5" heatid="22001" comment="aufgegeben nach 150m">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:02.74" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="288" birthdate="2006-01-01" gender="F" lastname="Hollatz" firstname="Ronja" license="0">
              <RESULTS>
                <RESULT resultid="888" eventid="11" swimtime="00:00:25.76" lane="1" heatid="11011" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="289" birthdate="2007-01-01" gender="F" lastname="Buse" firstname="Hermine" license="0">
              <RESULTS>
                <RESULT resultid="889" eventid="1" status="DSQ" swimtime="00:00:34.81" lane="5" heatid="1001" comment="Gesicht aus dem Wasser bei 35m" />
                <RESULT resultid="890" eventid="8" swimtime="00:01:15.69" lane="6" heatid="8008" />
                <RESULT resultid="891" eventid="11" swimtime="00:00:31.22" lane="2" heatid="11007" />
                <RESULT resultid="892" eventid="13" swimtime="00:02:52.36" lane="5" heatid="13005">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:16.69" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="893" eventid="16" swimtime="00:06:14.55" lane="1" heatid="16003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:22.67" />
                    <SPLIT distance="200" swimtime="00:03:00.39" />
                    <SPLIT distance="300" swimtime="00:04:39.31" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="894" eventid="18" swimtime="00:01:18.45" lane="7" heatid="18002" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="290" birthdate="2007-01-01" gender="M" lastname="Stuwe" firstname="Paul" license="0">
              <RESULTS>
                <RESULT resultid="895" eventid="2" swimtime="00:00:21.89" lane="6" heatid="2003" />
                <RESULT resultid="896" eventid="7" swimtime="00:09:18.37" lane="5" heatid="7002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:59.49" />
                    <SPLIT distance="200" swimtime="00:02:07.85" />
                    <SPLIT distance="300" swimtime="00:03:19.40" />
                    <SPLIT distance="400" swimtime="00:04:31.90" />
                    <SPLIT distance="500" swimtime="00:05:44.83" />
                    <SPLIT distance="600" swimtime="00:06:56.16" />
                    <SPLIT distance="700" swimtime="00:08:07.60" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="897" eventid="10" swimtime="00:04:29.70" lane="8" heatid="10002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:58.40" />
                    <SPLIT distance="200" swimtime="00:02:08.03" />
                    <SPLIT distance="300" swimtime="00:03:18.57" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="898" eventid="17" swimtime="00:04:40.70" lane="7" heatid="17003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:02.44" />
                    <SPLIT distance="200" swimtime="00:02:14.77" />
                    <SPLIT distance="300" swimtime="00:03:27.76" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="899" eventid="22" swimtime="00:18:27.07" lane="4" heatid="22001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:03.62" />
                    <SPLIT distance="200" swimtime="00:02:14.08" />
                    <SPLIT distance="300" swimtime="00:03:25.81" />
                    <SPLIT distance="400" swimtime="00:04:39.32" />
                    <SPLIT distance="500" swimtime="00:05:54.03" />
                    <SPLIT distance="600" swimtime="00:07:09.43" />
                    <SPLIT distance="700" swimtime="00:08:26.61" />
                    <SPLIT distance="800" swimtime="00:09:44.93" />
                    <SPLIT distance="900" swimtime="00:11:01.94" />
                    <SPLIT distance="1000" swimtime="00:12:16.84" />
                    <SPLIT distance="1100" swimtime="00:13:30.63" />
                    <SPLIT distance="1200" swimtime="00:14:46.64" />
                    <SPLIT distance="1300" swimtime="00:16:02.64" />
                    <SPLIT distance="1400" swimtime="00:17:15.58" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="291" birthdate="2008-01-01" gender="F" lastname="Liebhold" firstname="Lotta" license="0">
              <RESULTS>
                <RESULT resultid="900" eventid="1" swimtime="00:00:25.27" lane="2" heatid="1003" />
                <RESULT resultid="901" eventid="7" swimtime="00:10:37.77" lane="7" heatid="7002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:10.54" />
                    <SPLIT distance="200" swimtime="00:02:29.80" />
                    <SPLIT distance="300" swimtime="00:03:54.70" />
                    <SPLIT distance="400" swimtime="00:05:19.33" />
                    <SPLIT distance="500" swimtime="00:06:42.63" />
                    <SPLIT distance="600" swimtime="00:08:06.50" />
                    <SPLIT distance="700" swimtime="00:09:26.69" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="902" eventid="11" swimtime="00:00:26.52" lane="1" heatid="11010" />
                <RESULT resultid="903" eventid="16" swimtime="00:04:50.59" lane="3" heatid="16004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:08.23" />
                    <SPLIT distance="200" swimtime="00:02:23.92" />
                    <SPLIT distance="300" swimtime="00:03:40.64" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="904" eventid="18" swimtime="00:01:03.46" lane="2" heatid="18002" />
                <RESULT resultid="905" eventid="22" swimtime="00:21:01.32" lane="2" heatid="22001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:09.84" />
                    <SPLIT distance="200" swimtime="00:02:30.08" />
                    <SPLIT distance="300" swimtime="00:03:53.74" />
                    <SPLIT distance="400" swimtime="00:05:18.41" />
                    <SPLIT distance="500" swimtime="00:06:42.51" />
                    <SPLIT distance="600" swimtime="00:08:08.30" />
                    <SPLIT distance="700" swimtime="00:09:32.13" />
                    <SPLIT distance="800" swimtime="00:10:57.37" />
                    <SPLIT distance="900" swimtime="00:12:23.45" />
                    <SPLIT distance="1000" swimtime="00:13:52.04" />
                    <SPLIT distance="1100" swimtime="00:15:19.24" />
                    <SPLIT distance="1200" swimtime="00:16:51.05" />
                    <SPLIT distance="1300" swimtime="00:18:16.83" />
                    <SPLIT distance="1400" swimtime="00:19:42.01" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="292" birthdate="2009-01-01" gender="F" lastname="Weber" firstname="Augusta Swantje" license="0">
              <RESULTS>
                <RESULT resultid="906" eventid="1" status="DSQ" swimtime="00:00:28.67" lane="4" heatid="1001" comment="Gesicht aus dem Wasser bei 40m" />
                <RESULT resultid="907" eventid="8" swimtime="00:01:02.47" lane="8" heatid="8008" />
                <RESULT resultid="908" eventid="11" swimtime="00:00:27.95" lane="3" heatid="11008" />
                <RESULT resultid="909" eventid="13" swimtime="00:02:19.88" lane="5" heatid="13006">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:07.26" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="910" eventid="16" swimtime="00:05:10.98" lane="6" heatid="16003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:09.09" />
                    <SPLIT distance="200" swimtime="00:02:27.25" />
                    <SPLIT distance="300" swimtime="00:03:50.59" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="911" eventid="18" swimtime="00:01:10.04" lane="5" heatid="18001" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="294" birthdate="2010-01-01" gender="F" lastname="Rückert" firstname="Alma" license="0">
              <RESULTS>
                <RESULT resultid="913" eventid="3" swimtime="00:00:29.21" lane="7" heatid="3001" />
                <RESULT resultid="914" eventid="8" swimtime="00:01:06.82" lane="1" heatid="8007" />
                <RESULT resultid="915" eventid="11" swimtime="00:00:28.71" lane="1" heatid="11007" />
                <RESULT resultid="916" eventid="13" swimtime="00:02:32.45" lane="3" heatid="13005">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:13.16" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="917" eventid="16" swimtime="00:05:36.30" lane="4" heatid="16002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:15.42" />
                    <SPLIT distance="200" swimtime="00:02:45.39" />
                    <SPLIT distance="300" swimtime="00:04:16.72" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="918" eventid="18" swimtime="00:01:12.97" lane="2" heatid="18001" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="295" birthdate="2010-01-01" gender="F" lastname="Hoffmann" firstname="Lydia" license="0">
              <RESULTS>
                <RESULT resultid="919" eventid="3" swimtime="00:00:34.14" lane="1" heatid="3001" />
                <RESULT resultid="920" eventid="8" swimtime="00:01:16.36" lane="7" heatid="8006" />
                <RESULT resultid="921" eventid="11" swimtime="00:00:32.60" lane="7" heatid="11006" />
                <RESULT resultid="922" eventid="13" swimtime="00:02:50.82" lane="6" heatid="13004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:18.23" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="923" eventid="16" swimtime="00:05:53.63" lane="2" heatid="16002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:18.37" />
                    <SPLIT distance="200" swimtime="00:02:52.51" />
                    <SPLIT distance="300" swimtime="00:04:28.62" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="924" eventid="18" swimtime="00:01:20.06" lane="7" heatid="18001" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="296" birthdate="2010-01-01" gender="F" lastname="Schubert" firstname="Svea" license="0">
              <RESULTS>
                <RESULT resultid="925" eventid="3" swimtime="00:00:33.10" lane="8" heatid="3001" />
                <RESULT resultid="926" eventid="8" swimtime="00:01:09.52" lane="6" heatid="8006" />
                <RESULT resultid="927" eventid="11" swimtime="00:00:30.46" lane="5" heatid="11006" />
                <RESULT resultid="928" eventid="13" swimtime="00:02:35.59" lane="7" heatid="13005">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:16.07" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="929" eventid="16" swimtime="00:05:35.62" lane="8" heatid="16003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:20.10" />
                    <SPLIT distance="200" swimtime="00:02:47.81" />
                    <SPLIT distance="300" swimtime="00:04:13.17" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="930" eventid="18" swimtime="00:01:23.68" lane="8" heatid="18001" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="297" birthdate="2011-01-01" gender="M" lastname="Bartels" firstname="Constantin" license="0">
              <RESULTS>
                <RESULT resultid="931" eventid="9" swimtime="00:01:25.16" lane="6" heatid="9002" />
                <RESULT resultid="932" eventid="12" swimtime="00:00:38.16" lane="5" heatid="12001" />
                <RESULT resultid="933" eventid="14" swimtime="00:03:08.33" lane="2" heatid="14001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:29.91" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="934" eventid="17" swimtime="00:06:33.95" lane="3" heatid="17001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:29.05" />
                    <SPLIT distance="200" swimtime="00:03:10.86" />
                    <SPLIT distance="300" swimtime="00:04:52.60" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="298" birthdate="2011-01-01" gender="F" lastname="Wirsching" firstname="Ellen" license="0">
              <RESULTS>
                <RESULT resultid="935" eventid="8" swimtime="00:01:20.69" lane="3" heatid="8005" />
                <RESULT resultid="936" eventid="11" swimtime="00:00:34.59" lane="7" heatid="11005" />
                <RESULT resultid="937" eventid="13" swimtime="00:03:08.14" lane="3" heatid="13002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:28.10" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="938" eventid="16" swimtime="00:06:30.89" lane="3" heatid="16001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:28.05" />
                    <SPLIT distance="200" swimtime="00:03:08.59" />
                    <SPLIT distance="300" swimtime="00:04:51.64" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="299" birthdate="2011-01-01" gender="M" lastname="Knöfel" firstname="Florian" license="0">
              <RESULTS>
                <RESULT resultid="939" eventid="4" swimtime="00:00:34.32" lane="3" heatid="4001" />
                <RESULT resultid="940" eventid="9" swimtime="00:01:15.91" lane="2" heatid="9004" />
                <RESULT resultid="941" eventid="12" swimtime="00:00:32.79" lane="6" heatid="12003" />
                <RESULT resultid="942" eventid="14" swimtime="00:03:03.21" lane="4" heatid="14002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:28.27" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="943" eventid="17" swimtime="00:06:24.19" lane="7" heatid="17002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:27.33" />
                    <SPLIT distance="200" swimtime="00:03:06.46" />
                    <SPLIT distance="300" swimtime="00:04:45.33" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="944" eventid="19" swimtime="00:01:22.66" lane="3" heatid="19001" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="302" birthdate="2012-01-01" gender="F" lastname="Uhlig" firstname="Maike" license="0">
              <RESULTS>
                <RESULT resultid="947" eventid="5" swimtime="00:00:33.10" lane="7" heatid="5003" />
                <RESULT resultid="948" eventid="8" swimtime="00:01:16.21" lane="4" heatid="8003" />
                <RESULT resultid="949" eventid="11" swimtime="00:00:33.98" lane="2" heatid="11005" />
                <RESULT resultid="950" eventid="13" swimtime="00:02:57.82" lane="2" heatid="13003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:25.03" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="951" eventid="16" swimtime="00:06:25.73" lane="7" heatid="16002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:27.04" />
                    <SPLIT distance="200" swimtime="00:03:07.62" />
                    <SPLIT distance="300" swimtime="00:04:49.11" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="303" birthdate="2014-01-01" gender="F" lastname="Uhlig" firstname="Anna" license="0">
              <RESULTS>
                <RESULT resultid="952" eventid="5" swimtime="00:00:47.95" lane="7" heatid="5001" />
                <RESULT resultid="953" eventid="8" swimtime="00:01:34.74" lane="7" heatid="8001" />
                <RESULT resultid="954" eventid="11" swimtime="00:00:42.72" lane="7" heatid="11001" />
                <RESULT resultid="961" eventid="13" swimtime="00:03:34.51" lane="7" heatid="13002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:37.92" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY number="1" gender="M" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="874" eventid="21" swimtime="00:03:11.26" lane="1" heatid="21002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:55.92" />
                    <SPLIT distance="200" swimtime="00:01:45.25" />
                    <SPLIT distance="300" swimtime="00:02:29.41" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="290" number="1" />
                    <RELAYPOSITION athleteid="285" number="2" />
                    <RELAYPOSITION athleteid="287" number="3" />
                    <RELAYPOSITION athleteid="286" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" gender="F" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="912" eventid="20" swimtime="00:04:36.01" lane="2" heatid="20002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:09.69" />
                    <SPLIT distance="200" swimtime="00:02:17.90" />
                    <SPLIT distance="300" swimtime="00:03:32.87" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="296" number="1" />
                    <RELAYPOSITION athleteid="294" number="2" />
                    <RELAYPOSITION athleteid="295" number="3" />
                    <RELAYPOSITION athleteid="292" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
      </CLUBS>
    </MEET>
  </MEETS>
</LENEX>
