<?xml version="1.0" encoding="UTF-8"?>
<LENEX version="3.0">
  <CONSTRUCTOR name="EasyWk" version="5.23 BETA" registration="">
    <CONTACT name="Bjoern Stickan" internet="http://www.easywk.de" email="info@easywk.de" />
  </CONSTRUCTOR>
  <MEETS>
    <MEET city="Leipzig" course="LCM" name="63. Dt. Meisterschaften, 53. Dt. Jugendmeisterschaften, 44. Dt. Juniorenmeisterschaften, 11. Dt. Mastersmeisterschaften im Finswimming" nation="GER" organizer="SC DHfK Leipzig e.V., Abteilung Finswimming" hostclub="Verband Deutscher Sporttaucher e.V." deadline="2023-05-03" timing="AUTOMATIC">
      <CONTACT city="Leipzig" email="dm2023@egd-tb.de" fax="+49-341-4426911" name="Brandenburg, Thilo" phone="+49-178-8150839" street="Zum Leutzscher Holz 26" zip="04178" />
      <AGEDATE type="YEAR" value="2023-01-01" />
      <SESSIONS>
        <SESSION number="1" date="2023-05-12" daytime="13:55" officialmeeting="13:10" warmupfrom="12:15">
          <EVENTS>
            <EVENT eventid="1" number="1" gender="F" round="PRE">
              <SWIMSTYLE stroke="SURFACE" relaycount="1" distance="50" />
              <FEE value="650" currency="EUR" />
              <HEATS>
                <HEAT heatid="1001" number="1" />
                <HEAT heatid="1002" number="2" />
                <HEAT heatid="1003" number="3" />
                <HEAT heatid="1004" number="4" />
                <HEAT heatid="1005" number="5" />
                <HEAT heatid="1006" number="6" />
                <HEAT heatid="1007" number="7" />
                <HEAT heatid="1008" number="8" />
                <HEAT heatid="1009" number="9" />
                <HEAT heatid="1010" number="10" />
                <HEAT heatid="1011" number="11" />
                <HEAT heatid="1012" number="12" />
                <HEAT heatid="1013" number="13" />
                <HEAT heatid="1014" number="14" />
                <HEAT heatid="1015" number="15" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="4" agemax="13" agemin="12" name="Kategorie D">
                  <RANKINGS>
                    <RANKING place="9" resultid="234" />
                    <RANKING place="5" resultid="239" />
                    <RANKING place="18" resultid="303" />
                    <RANKING place="6" resultid="360" />
                    <RANKING place="11" resultid="371" />
                    <RANKING place="19" resultid="392" />
                    <RANKING place="4" resultid="492" />
                    <RANKING place="23" resultid="550" />
                    <RANKING place="2" resultid="570" />
                    <RANKING place="17" resultid="668" />
                    <RANKING place="14" resultid="698" />
                    <RANKING place="22" resultid="707" />
                    <RANKING place="7" resultid="725" />
                    <RANKING place="21" resultid="787" />
                    <RANKING place="15" resultid="791" />
                    <RANKING place="1" resultid="821" />
                    <RANKING place="13" resultid="832" />
                    <RANKING place="3" resultid="871" />
                    <RANKING place="10" resultid="877" />
                    <RANKING place="20" resultid="943" />
                    <RANKING place="8" resultid="1073" />
                    <RANKING place="26" resultid="1238" />
                    <RANKING place="27" resultid="1242" />
                    <RANKING place="12" resultid="1272" />
                    <RANKING place="25" resultid="1287" />
                    <RANKING place="16" resultid="1294" />
                    <RANKING place="24" resultid="1311" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3" agemax="15" agemin="14" name="Kategorie C">
                  <RANKINGS>
                    <RANKING place="17" resultid="153" />
                    <RANKING place="27" resultid="222" />
                    <RANKING place="11" resultid="273" />
                    <RANKING place="7" resultid="280" />
                    <RANKING place="12" resultid="284" />
                    <RANKING place="16" resultid="311" />
                    <RANKING place="6" resultid="376" />
                    <RANKING place="20" resultid="411" />
                    <RANKING place="14" resultid="437" />
                    <RANKING place="4" resultid="464" />
                    <RANKING place="18" resultid="488" />
                    <RANKING place="8" resultid="585" />
                    <RANKING place="22" resultid="597" />
                    <RANKING place="13" resultid="638" />
                    <RANKING place="25" resultid="841" />
                    <RANKING place="2" resultid="952" />
                    <RANKING place="3" resultid="1028" />
                    <RANKING place="10" resultid="1205" />
                    <RANKING place="5" resultid="1210" />
                    <RANKING place="1" resultid="1229" />
                    <RANKING place="24" resultid="1235" />
                    <RANKING place="26" resultid="1249" />
                    <RANKING place="9" resultid="1267" />
                    <RANKING place="21" resultid="1276" />
                    <RANKING place="15" resultid="1282" />
                    <RANKING place="28" resultid="1314" />
                    <RANKING place="23" resultid="1355" />
                    <RANKING place="19" resultid="1363" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2" agemax="17" agemin="16" name="Kategorie B">
                  <RANKINGS>
                    <RANKING place="12" resultid="50" />
                    <RANKING place="3" resultid="424" />
                    <RANKING place="15" resultid="433" />
                    <RANKING place="1" resultid="441" />
                    <RANKING place="14" resultid="517" />
                    <RANKING place="9" resultid="896" />
                    <RANKING place="16" resultid="956" />
                    <RANKING place="4" resultid="1049" />
                    <RANKING place="17" resultid="1095" />
                    <RANKING place="5" resultid="1096" />
                    <RANKING place="7" resultid="1137" />
                    <RANKING place="8" resultid="1147" />
                    <RANKING place="18" resultid="1151" />
                    <RANKING place="6" resultid="1163" />
                    <RANKING place="10" resultid="1191" />
                    <RANKING place="13" resultid="1224" />
                    <RANKING place="11" resultid="1318" />
                    <RANKING place="2" resultid="1342" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1" agemax="21" agemin="18" name="Junior:innen">
                  <RANKINGS>
                    <RANKING place="11" resultid="75" />
                    <RANKING place="16" resultid="106" />
                    <RANKING place="4" resultid="244" />
                    <RANKING place="10" resultid="255" />
                    <RANKING place="12" resultid="293" />
                    <RANKING place="13" resultid="454" />
                    <RANKING place="8" resultid="534" />
                    <RANKING place="6" resultid="744" />
                    <RANKING place="3" resultid="758" />
                    <RANKING place="9" resultid="765" />
                    <RANKING place="14" resultid="853" />
                    <RANKING place="7" resultid="864" />
                    <RANKING place="15" resultid="882" />
                    <RANKING place="2" resultid="974" />
                    <RANKING place="16" resultid="1033" />
                    <RANKING place="4" resultid="1126" />
                    <RANKING place="1" resultid="1143" />
                    <RANKING place="18" resultid="1180" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="34" agemin="29" name="Master A">
                  <RANKINGS>
                    <RANKING place="1" resultid="3" />
                    <RANKING place="2" resultid="46" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6" agemax="44" agemin="35" name="Master B">
                  <RANKINGS>
                    <RANKING place="2" resultid="647" />
                    <RANKING place="3" resultid="653" />
                    <RANKING place="4" resultid="772" />
                    <RANKING place="1" resultid="996" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7" agemax="54" agemin="45" name="Master C">
                  <RANKINGS>
                    <RANKING place="2" resultid="26" />
                    <RANKING place="3" resultid="836" />
                    <RANKING place="1" resultid="1019" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8" agemax="64" agemin="55" name="Master D">
                  <RANKINGS>
                    <RANKING place="1" resultid="657" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9" agemax="-1" agemin="65" name="Master E">
                  <RANKINGS>
                    <RANKING place="1" resultid="992" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10" agemax="-1" agemin="12" name="offene Wertung">
                  <RANKINGS>
                    <RANKING place="40" resultid="3" />
                    <RANKING place="66" resultid="26" />
                    <RANKING place="93" resultid="46" />
                    <RANKING place="43" resultid="50" />
                    <RANKING place="23" resultid="75" />
                    <RANKING place="26" resultid="82" />
                    <RANKING place="43" resultid="106" />
                    <RANKING place="64" resultid="153" />
                    <RANKING place="95" resultid="222" />
                    <RANKING place="73" resultid="234" />
                    <RANKING place="65" resultid="239" />
                    <RANKING place="6" resultid="244" />
                    <RANKING place="21" resultid="255" />
                    <RANKING place="50" resultid="273" />
                    <RANKING place="30" resultid="280" />
                    <RANKING place="52" resultid="284" />
                    <RANKING place="41" resultid="288" />
                    <RANKING place="27" resultid="293" />
                    <RANKING place="94" resultid="303" />
                    <RANKING place="62" resultid="311" />
                    <RANKING place="68" resultid="360" />
                    <RANKING place="77" resultid="371" />
                    <RANKING place="28" resultid="376" />
                    <RANKING place="97" resultid="392" />
                    <RANKING place="76" resultid="411" />
                    <RANKING place="11" resultid="424" />
                    <RANKING place="51" resultid="433" />
                    <RANKING place="57" resultid="437" />
                    <RANKING place="8" resultid="441" />
                    <RANKING place="31" resultid="454" />
                    <RANKING place="22" resultid="464" />
                    <RANKING place="72" resultid="488" />
                    <RANKING place="63" resultid="492" />
                    <RANKING place="49" resultid="517" />
                    <RANKING place="16" resultid="534" />
                    <RANKING place="101" resultid="550" />
                    <RANKING place="47" resultid="570" />
                    <RANKING place="36" resultid="585" />
                    <RANKING place="83" resultid="597" />
                    <RANKING place="55" resultid="638" />
                    <RANKING place="67" resultid="647" />
                    <RANKING place="90" resultid="653" />
                    <RANKING place="106" resultid="657" />
                    <RANKING place="89" resultid="668" />
                    <RANKING place="82" resultid="698" />
                    <RANKING place="100" resultid="707" />
                    <RANKING place="69" resultid="725" />
                    <RANKING place="10" resultid="744" />
                    <RANKING place="5" resultid="758" />
                    <RANKING place="19" resultid="765" />
                    <RANKING place="92" resultid="772" />
                    <RANKING place="4" resultid="777" />
                    <RANKING place="99" resultid="787" />
                    <RANKING place="84" resultid="791" />
                    <RANKING place="46" resultid="821" />
                    <RANKING place="81" resultid="832" />
                    <RANKING place="70" resultid="836" />
                    <RANKING place="88" resultid="841" />
                    <RANKING place="33" resultid="853" />
                    <RANKING place="14" resultid="864" />
                    <RANKING place="53" resultid="871" />
                    <RANKING place="75" resultid="877" />
                    <RANKING place="39" resultid="882" />
                    <RANKING place="32" resultid="896" />
                    <RANKING place="33" resultid="927" />
                    <RANKING place="98" resultid="943" />
                    <RANKING place="17" resultid="950" />
                    <RANKING place="18" resultid="952" />
                    <RANKING place="56" resultid="956" />
                    <RANKING place="2" resultid="974" />
                    <RANKING place="105" resultid="992" />
                    <RANKING place="61" resultid="996" />
                    <RANKING place="59" resultid="1019" />
                    <RANKING place="20" resultid="1028" />
                    <RANKING place="43" resultid="1033" />
                    <RANKING place="12" resultid="1049" />
                    <RANKING place="71" resultid="1073" />
                    <RANKING place="60" resultid="1095" />
                    <RANKING place="13" resultid="1096" />
                    <RANKING place="6" resultid="1126" />
                    <RANKING place="24" resultid="1137" />
                    <RANKING place="1" resultid="1143" />
                    <RANKING place="29" resultid="1147" />
                    <RANKING place="80" resultid="1151" />
                    <RANKING place="15" resultid="1163" />
                    <RANKING place="54" resultid="1180" />
                    <RANKING place="35" resultid="1191" />
                    <RANKING place="42" resultid="1205" />
                    <RANKING place="25" resultid="1210" />
                    <RANKING place="48" resultid="1224" />
                    <RANKING place="3" resultid="1229" />
                    <RANKING place="87" resultid="1235" />
                    <RANKING place="104" resultid="1238" />
                    <RANKING place="107" resultid="1242" />
                    <RANKING place="91" resultid="1249" />
                    <RANKING place="38" resultid="1267" />
                    <RANKING place="78" resultid="1272" />
                    <RANKING place="79" resultid="1276" />
                    <RANKING place="58" resultid="1282" />
                    <RANKING place="103" resultid="1287" />
                    <RANKING place="85" resultid="1294" />
                    <RANKING place="102" resultid="1311" />
                    <RANKING place="96" resultid="1314" />
                    <RANKING place="37" resultid="1318" />
                    <RANKING place="9" resultid="1342" />
                    <RANKING place="86" resultid="1355" />
                    <RANKING place="74" resultid="1363" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11" agemax="-1" agemin="12" name="Internationale offene Wertung">
                  <RANKINGS>
                    <RANKING place="44" resultid="3" />
                    <RANKING place="73" resultid="26" />
                    <RANKING place="53" resultid="39" />
                    <RANKING place="101" resultid="46" />
                    <RANKING place="47" resultid="50" />
                    <RANKING place="25" resultid="75" />
                    <RANKING place="28" resultid="82" />
                    <RANKING place="47" resultid="106" />
                    <RANKING place="69" resultid="153" />
                    <RANKING place="30" resultid="171" />
                    <RANKING place="77" resultid="213" />
                    <RANKING place="103" resultid="222" />
                    <RANKING place="81" resultid="234" />
                    <RANKING place="70" resultid="239" />
                    <RANKING place="7" resultid="244" />
                    <RANKING place="23" resultid="255" />
                    <RANKING place="55" resultid="273" />
                    <RANKING place="33" resultid="280" />
                    <RANKING place="57" resultid="284" />
                    <RANKING place="45" resultid="288" />
                    <RANKING place="29" resultid="293" />
                    <RANKING place="102" resultid="303" />
                    <RANKING place="67" resultid="311" />
                    <RANKING place="75" resultid="360" />
                    <RANKING place="85" resultid="371" />
                    <RANKING place="31" resultid="376" />
                    <RANKING place="105" resultid="392" />
                    <RANKING place="84" resultid="411" />
                    <RANKING place="12" resultid="424" />
                    <RANKING place="56" resultid="433" />
                    <RANKING place="62" resultid="437" />
                    <RANKING place="9" resultid="441" />
                    <RANKING place="34" resultid="454" />
                    <RANKING place="72" resultid="459" />
                    <RANKING place="24" resultid="464" />
                    <RANKING place="80" resultid="488" />
                    <RANKING place="68" resultid="492" />
                    <RANKING place="53" resultid="517" />
                    <RANKING place="17" resultid="534" />
                    <RANKING place="109" resultid="550" />
                    <RANKING place="51" resultid="570" />
                    <RANKING place="40" resultid="575" />
                    <RANKING place="39" resultid="585" />
                    <RANKING place="91" resultid="597" />
                    <RANKING place="60" resultid="638" />
                    <RANKING place="74" resultid="647" />
                    <RANKING place="98" resultid="653" />
                    <RANKING place="114" resultid="657" />
                    <RANKING place="97" resultid="668" />
                    <RANKING place="90" resultid="698" />
                    <RANKING place="108" resultid="707" />
                    <RANKING place="76" resultid="725" />
                    <RANKING place="11" resultid="744" />
                    <RANKING place="6" resultid="758" />
                    <RANKING place="21" resultid="765" />
                    <RANKING place="100" resultid="772" />
                    <RANKING place="4" resultid="777" />
                    <RANKING place="107" resultid="787" />
                    <RANKING place="92" resultid="791" />
                    <RANKING place="50" resultid="821" />
                    <RANKING place="89" resultid="832" />
                    <RANKING place="78" resultid="836" />
                    <RANKING place="96" resultid="841" />
                    <RANKING place="36" resultid="853" />
                    <RANKING place="15" resultid="864" />
                    <RANKING place="58" resultid="871" />
                    <RANKING place="83" resultid="877" />
                    <RANKING place="43" resultid="882" />
                    <RANKING place="35" resultid="896" />
                    <RANKING place="36" resultid="927" />
                    <RANKING place="106" resultid="943" />
                    <RANKING place="19" resultid="950" />
                    <RANKING place="20" resultid="952" />
                    <RANKING place="61" resultid="956" />
                    <RANKING place="5" resultid="960" />
                    <RANKING place="2" resultid="974" />
                    <RANKING place="71" resultid="978" />
                    <RANKING place="113" resultid="992" />
                    <RANKING place="66" resultid="996" />
                    <RANKING place="64" resultid="1019" />
                    <RANKING place="22" resultid="1028" />
                    <RANKING place="47" resultid="1033" />
                    <RANKING place="13" resultid="1049" />
                    <RANKING place="79" resultid="1073" />
                    <RANKING place="65" resultid="1095" />
                    <RANKING place="14" resultid="1096" />
                    <RANKING place="7" resultid="1126" />
                    <RANKING place="26" resultid="1137" />
                    <RANKING place="1" resultid="1143" />
                    <RANKING place="32" resultid="1147" />
                    <RANKING place="88" resultid="1151" />
                    <RANKING place="18" resultid="1158" />
                    <RANKING place="16" resultid="1163" />
                    <RANKING place="59" resultid="1180" />
                    <RANKING place="38" resultid="1191" />
                    <RANKING place="46" resultid="1205" />
                    <RANKING place="27" resultid="1210" />
                    <RANKING place="52" resultid="1224" />
                    <RANKING place="3" resultid="1229" />
                    <RANKING place="95" resultid="1235" />
                    <RANKING place="112" resultid="1238" />
                    <RANKING place="115" resultid="1242" />
                    <RANKING place="99" resultid="1249" />
                    <RANKING place="42" resultid="1267" />
                    <RANKING place="86" resultid="1272" />
                    <RANKING place="87" resultid="1276" />
                    <RANKING place="63" resultid="1282" />
                    <RANKING place="111" resultid="1287" />
                    <RANKING place="93" resultid="1294" />
                    <RANKING place="110" resultid="1311" />
                    <RANKING place="104" resultid="1314" />
                    <RANKING place="41" resultid="1318" />
                    <RANKING place="10" resultid="1342" />
                    <RANKING place="94" resultid="1355" />
                    <RANKING place="82" resultid="1363" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="2" number="2" gender="M" round="PRE">
              <SWIMSTYLE stroke="SURFACE" relaycount="1" distance="50" />
              <FEE value="650" currency="EUR" />
              <HEATS>
                <HEAT heatid="2001" number="1" />
                <HEAT heatid="2002" number="2" />
                <HEAT heatid="2003" number="3" />
                <HEAT heatid="2004" number="4" />
                <HEAT heatid="2005" number="5" />
                <HEAT heatid="2006" number="6" />
                <HEAT heatid="2007" number="7" />
                <HEAT heatid="2008" number="8" />
                <HEAT heatid="2009" number="9" />
                <HEAT heatid="2010" number="10" />
                <HEAT heatid="2011" number="11" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="4" agemax="13" agemin="12" name="Kategorie D">
                  <RANKINGS>
                    <RANKING place="9" resultid="92" />
                    <RANKING place="6" resultid="266" />
                    <RANKING place="10" resultid="590" />
                    <RANKING place="1" resultid="613" />
                    <RANKING place="3" resultid="620" />
                    <RANKING place="11" resultid="630" />
                    <RANKING place="4" resultid="672" />
                    <RANKING place="2" resultid="701" />
                    <RANKING place="8" resultid="730" />
                    <RANKING place="7" resultid="1089" />
                    <RANKING place="12" resultid="1093" />
                    <RANKING place="16" resultid="1108" />
                    <RANKING place="13" resultid="1187" />
                    <RANKING place="15" resultid="1246" />
                    <RANKING place="14" resultid="1298" />
                    <RANKING place="5" resultid="1303" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3" agemax="15" agemin="14" name="Kategorie C">
                  <RANKINGS>
                    <RANKING place="16" resultid="112" />
                    <RANKING place="9" resultid="121" />
                    <RANKING place="14" resultid="126" />
                    <RANKING place="11" resultid="397" />
                    <RANKING place="4" resultid="415" />
                    <RANKING place="19" resultid="498" />
                    <RANKING place="7" resultid="506" />
                    <RANKING place="10" resultid="522" />
                    <RANKING place="2" resultid="527" />
                    <RANKING place="17" resultid="604" />
                    <RANKING place="15" resultid="681" />
                    <RANKING place="3" resultid="715" />
                    <RANKING place="13" resultid="848" />
                    <RANKING place="18" resultid="856" />
                    <RANKING place="5" resultid="915" />
                    <RANKING place="7" resultid="1105" />
                    <RANKING place="6" resultid="1196" />
                    <RANKING place="12" resultid="1216" />
                    <RANKING place="20" resultid="1290" />
                    <RANKING place="1" resultid="1350" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2" agemax="17" agemin="16" name="Kategorie B">
                  <RANKINGS>
                    <RANKING place="5" resultid="261" />
                    <RANKING place="2" resultid="633" />
                    <RANKING place="8" resultid="684" />
                    <RANKING place="6" resultid="720" />
                    <RANKING place="1" resultid="795" />
                    <RANKING place="3" resultid="922" />
                    <RANKING place="7" resultid="1081" />
                    <RANKING place="4" resultid="1117" />
                    <RANKING place="9" resultid="1368" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1" agemax="21" agemin="18" name="Junior:innen">
                  <RANKINGS>
                    <RANKING place="8" resultid="19" />
                    <RANKING place="10" resultid="187" />
                    <RANKING place="11" resultid="298" />
                    <RANKING place="12" resultid="307" />
                    <RANKING place="9" resultid="316" />
                    <RANKING place="1" resultid="386" />
                    <RANKING place="6" resultid="430" />
                    <RANKING place="2" resultid="474" />
                    <RANKING place="7" resultid="860" />
                    <RANKING place="5" resultid="1201" />
                    <RANKING place="4" resultid="1220" />
                    <RANKING place="3" resultid="1260" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="34" agemin="29" name="Master A">
                  <RANKINGS>
                    <RANKING place="1" resultid="965" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6" agemax="44" agemin="35" name="Master B">
                  <RANKINGS>
                    <RANKING place="3" resultid="32" />
                    <RANKING place="2" resultid="1092" />
                    <RANKING place="1" resultid="1382" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7" agemax="54" agemin="45" name="Master C">
                  <RANKINGS>
                    <RANKING place="4" resultid="179" />
                    <RANKING place="6" resultid="539" />
                    <RANKING place="5" resultid="608" />
                    <RANKING place="2" resultid="782" />
                    <RANKING place="3" resultid="891" />
                    <RANKING place="1" resultid="1008" />
                    <RANKING place="7" resultid="1014" />
                    <RANKING place="8" resultid="1375" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8" agemax="64" agemin="55" name="Master D">
                  <RANKINGS>
                    <RANKING place="1" resultid="9" />
                    <RANKING place="3" resultid="197" />
                    <RANKING place="4" resultid="479" />
                    <RANKING place="5" resultid="735" />
                    <RANKING place="6" resultid="827" />
                    <RANKING place="2" resultid="1024" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9" agemax="-1" agemin="65" name="Master E">
                  <RANKINGS>
                    <RANKING place="1" resultid="192" />
                    <RANKING place="2" resultid="750" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10" agemax="-1" agemin="12" name="offene Wertung">
                  <RANKINGS>
                    <RANKING place="30" resultid="9" />
                    <RANKING place="19" resultid="19" />
                    <RANKING place="48" resultid="32" />
                    <RANKING place="69" resultid="92" />
                    <RANKING place="62" resultid="112" />
                    <RANKING place="38" resultid="121" />
                    <RANKING place="58" resultid="126" />
                    <RANKING place="43" resultid="179" />
                    <RANKING place="24" resultid="187" />
                    <RANKING place="60" resultid="192" />
                    <RANKING place="45" resultid="197" />
                    <RANKING place="21" resultid="261" />
                    <RANKING place="64" resultid="266" />
                    <RANKING place="31" resultid="298" />
                    <RANKING place="44" resultid="307" />
                    <RANKING place="20" resultid="316" />
                    <RANKING place="5" resultid="386" />
                    <RANKING place="53" resultid="397" />
                    <RANKING place="25" resultid="415" />
                    <RANKING place="16" resultid="430" />
                    <RANKING place="9" resultid="474" />
                    <RANKING place="47" resultid="479" />
                    <RANKING place="70" resultid="498" />
                    <RANKING place="35" resultid="506" />
                    <RANKING place="42" resultid="522" />
                    <RANKING place="14" resultid="527" />
                    <RANKING place="49" resultid="539" />
                    <RANKING place="8" resultid="556" />
                    <RANKING place="72" resultid="590" />
                    <RANKING place="64" resultid="604" />
                    <RANKING place="46" resultid="608" />
                    <RANKING place="50" resultid="613" />
                    <RANKING place="56" resultid="620" />
                    <RANKING place="73" resultid="630" />
                    <RANKING place="3" resultid="633" />
                    <RANKING place="61" resultid="672" />
                    <RANKING place="59" resultid="681" />
                    <RANKING place="33" resultid="684" />
                    <RANKING place="51" resultid="701" />
                    <RANKING place="23" resultid="715" />
                    <RANKING place="26" resultid="720" />
                    <RANKING place="68" resultid="730" />
                    <RANKING place="71" resultid="735" />
                    <RANKING place="79" resultid="750" />
                    <RANKING place="37" resultid="782" />
                    <RANKING place="1" resultid="795" />
                    <RANKING place="74" resultid="827" />
                    <RANKING place="57" resultid="848" />
                    <RANKING place="67" resultid="856" />
                    <RANKING place="18" resultid="860" />
                    <RANKING place="16" resultid="887" />
                    <RANKING place="40" resultid="891" />
                    <RANKING place="27" resultid="915" />
                    <RANKING place="6" resultid="922" />
                    <RANKING place="7" resultid="939" />
                    <RANKING place="2" resultid="965" />
                    <RANKING place="4" resultid="987" />
                    <RANKING place="22" resultid="1008" />
                    <RANKING place="52" resultid="1014" />
                    <RANKING place="38" resultid="1024" />
                    <RANKING place="28" resultid="1081" />
                    <RANKING place="66" resultid="1089" />
                    <RANKING place="34" resultid="1092" />
                    <RANKING place="75" resultid="1093" />
                    <RANKING place="35" resultid="1105" />
                    <RANKING place="81" resultid="1108" />
                    <RANKING place="13" resultid="1117" />
                    <RANKING place="76" resultid="1187" />
                    <RANKING place="32" resultid="1196" />
                    <RANKING place="15" resultid="1201" />
                    <RANKING place="54" resultid="1216" />
                    <RANKING place="12" resultid="1220" />
                    <RANKING place="80" resultid="1246" />
                    <RANKING place="10" resultid="1260" />
                    <RANKING place="77" resultid="1290" />
                    <RANKING place="78" resultid="1298" />
                    <RANKING place="62" resultid="1303" />
                    <RANKING place="11" resultid="1350" />
                    <RANKING place="41" resultid="1368" />
                    <RANKING place="54" resultid="1375" />
                    <RANKING place="29" resultid="1382" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11" agemax="-1" agemin="12" name="Internationale offene Wertung">
                  <RANKINGS>
                    <RANKING place="32" resultid="9" />
                    <RANKING place="21" resultid="19" />
                    <RANKING place="50" resultid="32" />
                    <RANKING place="71" resultid="92" />
                    <RANKING place="64" resultid="112" />
                    <RANKING place="40" resultid="121" />
                    <RANKING place="60" resultid="126" />
                    <RANKING place="45" resultid="179" />
                    <RANKING place="26" resultid="187" />
                    <RANKING place="62" resultid="192" />
                    <RANKING place="47" resultid="197" />
                    <RANKING place="23" resultid="261" />
                    <RANKING place="66" resultid="266" />
                    <RANKING place="33" resultid="298" />
                    <RANKING place="46" resultid="307" />
                    <RANKING place="22" resultid="316" />
                    <RANKING place="5" resultid="386" />
                    <RANKING place="55" resultid="397" />
                    <RANKING place="27" resultid="415" />
                    <RANKING place="18" resultid="430" />
                    <RANKING place="9" resultid="474" />
                    <RANKING place="49" resultid="479" />
                    <RANKING place="72" resultid="498" />
                    <RANKING place="37" resultid="506" />
                    <RANKING place="44" resultid="522" />
                    <RANKING place="16" resultid="527" />
                    <RANKING place="51" resultid="539" />
                    <RANKING place="8" resultid="556" />
                    <RANKING place="74" resultid="590" />
                    <RANKING place="66" resultid="604" />
                    <RANKING place="48" resultid="608" />
                    <RANKING place="52" resultid="613" />
                    <RANKING place="58" resultid="620" />
                    <RANKING place="75" resultid="630" />
                    <RANKING place="3" resultid="633" />
                    <RANKING place="63" resultid="672" />
                    <RANKING place="61" resultid="681" />
                    <RANKING place="35" resultid="684" />
                    <RANKING place="53" resultid="701" />
                    <RANKING place="25" resultid="715" />
                    <RANKING place="28" resultid="720" />
                    <RANKING place="70" resultid="730" />
                    <RANKING place="73" resultid="735" />
                    <RANKING place="81" resultid="750" />
                    <RANKING place="39" resultid="782" />
                    <RANKING place="1" resultid="795" />
                    <RANKING place="76" resultid="827" />
                    <RANKING place="59" resultid="848" />
                    <RANKING place="69" resultid="856" />
                    <RANKING place="20" resultid="860" />
                    <RANKING place="18" resultid="887" />
                    <RANKING place="42" resultid="891" />
                    <RANKING place="29" resultid="915" />
                    <RANKING place="6" resultid="922" />
                    <RANKING place="7" resultid="939" />
                    <RANKING place="2" resultid="965" />
                    <RANKING place="15" resultid="970" />
                    <RANKING place="4" resultid="987" />
                    <RANKING place="24" resultid="1008" />
                    <RANKING place="54" resultid="1014" />
                    <RANKING place="40" resultid="1024" />
                    <RANKING place="30" resultid="1081" />
                    <RANKING place="68" resultid="1089" />
                    <RANKING place="36" resultid="1092" />
                    <RANKING place="77" resultid="1093" />
                    <RANKING place="37" resultid="1105" />
                    <RANKING place="83" resultid="1108" />
                    <RANKING place="13" resultid="1117" />
                    <RANKING place="13" resultid="1170" />
                    <RANKING place="78" resultid="1187" />
                    <RANKING place="34" resultid="1196" />
                    <RANKING place="17" resultid="1201" />
                    <RANKING place="56" resultid="1216" />
                    <RANKING place="12" resultid="1220" />
                    <RANKING place="82" resultid="1246" />
                    <RANKING place="10" resultid="1260" />
                    <RANKING place="79" resultid="1290" />
                    <RANKING place="80" resultid="1298" />
                    <RANKING place="64" resultid="1303" />
                    <RANKING place="11" resultid="1350" />
                    <RANKING place="43" resultid="1368" />
                    <RANKING place="56" resultid="1375" />
                    <RANKING place="31" resultid="1382" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="3" number="3" gender="F" round="TIM">
              <SWIMSTYLE stroke="SURFACE" relaycount="1" distance="1500" />
              <FEE value="650" currency="EUR" />
              <HEATS>
                <HEAT heatid="3001" number="1" />
                <HEAT heatid="3002" number="2" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="4" agemax="13" agemin="12" name="Kategorie D">
                  <RANKINGS>
                    <RANKING place="2" resultid="420" />
                    <RANKING place="3" resultid="545" />
                    <RANKING place="1" resultid="822" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3" agemax="15" agemin="14" name="Kategorie C">
                  <RANKINGS>
                    <RANKING place="1" resultid="639" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2" agemax="17" agemin="16" name="Kategorie B">
                  <RANKINGS>
                    <RANKING place="2" resultid="51" />
                    <RANKING place="5" resultid="381" />
                    <RANKING place="4" resultid="1100" />
                    <RANKING place="3" resultid="1138" />
                    <RANKING place="1" resultid="1164" />
                    <RANKING place="6" resultid="1253" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1" agemax="21" agemin="18" name="Junior:innen">
                  <RANKINGS>
                    <RANKING place="1" resultid="147" />
                    <RANKING place="2" resultid="1060" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10" agemax="-1" agemin="12" name="offene Wertung">
                  <RANKINGS>
                    <RANKING place="4" resultid="51" />
                    <RANKING place="2" resultid="116" />
                    <RANKING place="7" resultid="140" />
                    <RANKING place="3" resultid="147" />
                    <RANKING place="8" resultid="381" />
                    <RANKING place="13" resultid="420" />
                    <RANKING place="14" resultid="545" />
                    <RANKING place="11" resultid="639" />
                    <RANKING place="12" resultid="822" />
                    <RANKING place="10" resultid="1060" />
                    <RANKING place="6" resultid="1100" />
                    <RANKING place="5" resultid="1138" />
                    <RANKING place="1" resultid="1164" />
                    <RANKING place="9" resultid="1253" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11" agemax="-1" agemin="12" name="Internationale offene Wertung">
                  <RANKINGS>
                    <RANKING place="4" resultid="51" />
                    <RANKING place="2" resultid="116" />
                    <RANKING place="7" resultid="140" />
                    <RANKING place="3" resultid="147" />
                    <RANKING place="8" resultid="381" />
                    <RANKING place="13" resultid="420" />
                    <RANKING place="14" resultid="545" />
                    <RANKING place="11" resultid="639" />
                    <RANKING place="12" resultid="822" />
                    <RANKING place="10" resultid="1060" />
                    <RANKING place="6" resultid="1100" />
                    <RANKING place="5" resultid="1138" />
                    <RANKING place="1" resultid="1164" />
                    <RANKING place="9" resultid="1253" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="4" number="4" gender="M" round="TIM">
              <SWIMSTYLE stroke="SURFACE" relaycount="1" distance="1500" />
              <FEE value="650" currency="EUR" />
              <HEATS>
                <HEAT heatid="4001" number="1" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="4" agemax="13" agemin="12" name="Kategorie D">
                  <RANKINGS>
                    <RANKING place="1" resultid="93" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3" agemax="15" agemin="14" name="Kategorie C">
                  <RANKINGS>
                    <RANKING place="2" resultid="127" />
                    <RANKING place="1" resultid="448" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2" agemax="17" agemin="16" name="Kategorie B">
                  <RANKINGS>
                    <RANKING place="1" resultid="1369" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1" agemax="21" agemin="18" name="Junior:innen" />
                <AGEGROUP agegroupid="10" agemax="-1" agemin="12" name="offene Wertung">
                  <RANKINGS>
                    <RANKING place="4" resultid="93" />
                    <RANKING place="2" resultid="127" />
                    <RANKING place="1" resultid="448" />
                    <RANKING place="3" resultid="1369" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="5" number="201" gender="F" round="TIM">
              <SWIMSTYLE stroke="BIFIN" relaycount="1" distance="100" />
              <FEE value="1000" currency="EUR" />
              <HEATS>
                <HEAT heatid="5001" number="1" />
                <HEAT heatid="5002" number="2" />
                <HEAT heatid="5003" number="3" />
                <HEAT heatid="5004" number="4" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="-1" agemin="12" name="offene Klasse">
                  <RANKINGS>
                    <RANKING place="3" resultid="80" />
                    <RANKING place="2" resultid="87" />
                    <RANKING place="18" resultid="216" />
                    <RANKING place="23" resultid="395" />
                    <RANKING place="9" resultid="457" />
                    <RANKING place="13" resultid="462" />
                    <RANKING place="19" resultid="497" />
                    <RANKING place="25" resultid="554" />
                    <RANKING place="7" resultid="581" />
                    <RANKING place="16" resultid="583" />
                    <RANKING place="15" resultid="655" />
                    <RANKING place="21" resultid="662" />
                    <RANKING place="1" resultid="763" />
                    <RANKING place="12" resultid="847" />
                    <RANKING place="5" resultid="855" />
                    <RANKING place="6" resultid="875" />
                    <RANKING place="10" resultid="886" />
                    <RANKING place="8" resultid="903" />
                    <RANKING place="24" resultid="994" />
                    <RANKING place="17" resultid="998" />
                    <RANKING place="14" resultid="1022" />
                    <RANKING place="4" resultid="1214" />
                    <RANKING place="20" resultid="1240" />
                    <RANKING place="22" resultid="1313" />
                    <RANKING place="11" resultid="1378" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="6" number="202" gender="M" round="TIM">
              <SWIMSTYLE stroke="BIFIN" relaycount="1" distance="100" />
              <FEE value="1000" currency="EUR" />
              <HEATS>
                <HEAT heatid="6001" number="1" />
                <HEAT heatid="6002" number="2" />
                <HEAT heatid="6003" number="3" />
                <HEAT heatid="6004" number="4" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="-1" agemin="12" name="offene Klasse">
                  <RANKINGS>
                    <RANKING place="12" resultid="17" />
                    <RANKING place="10" resultid="37" />
                    <RANKING place="18" resultid="105" />
                    <RANKING place="2" resultid="165" />
                    <RANKING place="3" resultid="169" />
                    <RANKING place="21" resultid="185" />
                    <RANKING place="5" resultid="190" />
                    <RANKING place="19" resultid="206" />
                    <RANKING place="7" resultid="211" />
                    <RANKING place="4" resultid="220" />
                    <RANKING place="11" resultid="482" />
                    <RANKING place="23" resultid="500" />
                    <RANKING place="13" resultid="512" />
                    <RANKING place="16" resultid="543" />
                    <RANKING place="1" resultid="560" />
                    <RANKING place="8" resultid="688" />
                    <RANKING place="25" resultid="736" />
                    <RANKING place="6" resultid="785" />
                    <RANKING place="26" resultid="831" />
                    <RANKING place="24" resultid="858" />
                    <RANKING place="17" resultid="1002" />
                    <RANKING place="20" resultid="1006" />
                    <RANKING place="9" resultid="1012" />
                    <RANKING place="22" resultid="1017" />
                    <RANKING place="15" resultid="1026" />
                    <RANKING place="14" resultid="1379" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="7" number="101" gender="F" round="FIN">
              <SWIMSTYLE stroke="SURFACE" relaycount="1" distance="50" />
              <HEATS>
                <HEAT heatid="7001" number="1" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="10" agemax="-1" agemin="12" name="offene Wertung">
                  <RANKINGS>
                    <RANKING place="2" resultid="1404" />
                    <RANKING place="3" resultid="1405" />
                    <RANKING place="1" resultid="1407" />
                    <RANKING place="6" resultid="1409" />
                    <RANKING place="5" resultid="1410" />
                    <RANKING place="4" resultid="1411" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11" agemax="-1" agemin="12" name="Internationale offene Wertung">
                  <RANKINGS>
                    <RANKING place="2" resultid="1404" />
                    <RANKING place="4" resultid="1405" />
                    <RANKING place="1" resultid="1407" />
                    <RANKING place="2" resultid="1408" />
                    <RANKING place="7" resultid="1409" />
                    <RANKING place="6" resultid="1410" />
                    <RANKING place="5" resultid="1411" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="8" number="102" gender="M" round="FIN">
              <SWIMSTYLE stroke="SURFACE" relaycount="1" distance="50" />
              <HEATS>
                <HEAT heatid="8001" number="1" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="10" agemax="-1" agemin="12" name="offene Wertung">
                  <RANKINGS>
                    <RANKING place="2" resultid="1412" />
                    <RANKING place="1" resultid="1413" />
                    <RANKING place="3" resultid="1414" />
                    <RANKING place="4" resultid="1415" />
                    <RANKING place="5" resultid="1416" />
                    <RANKING place="7" resultid="1417" />
                    <RANKING place="6" resultid="1418" />
                    <RANKING place="8" resultid="1419" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="9" number="303" gender="F" round="FIN">
              <SWIMSTYLE stroke="SURFACE" relaycount="1" distance="1500" />
              <FEE value="650" currency="EUR" />
              <HEATS>
                <HEAT heatid="9001" number="1" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="4" agemax="13" agemin="12" name="Kategorie D" />
                <AGEGROUP agegroupid="3" agemax="15" agemin="14" name="Kategorie C" />
                <AGEGROUP agegroupid="2" agemax="17" agemin="16" name="Kategorie B">
                  <RANKINGS>
                    <RANKING place="2" resultid="228" />
                    <RANKING place="1" resultid="934" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1" agemax="21" agemin="18" name="Junior:innen">
                  <RANKINGS>
                    <RANKING place="3" resultid="107" />
                    <RANKING place="2" resultid="1127" />
                    <RANKING place="1" resultid="1132" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10" agemax="-1" agemin="12" name="offene Wertung">
                  <RANKINGS>
                    <RANKING place="3" resultid="59" />
                    <RANKING place="6" resultid="107" />
                    <RANKING place="4" resultid="228" />
                    <RANKING place="2" resultid="934" />
                    <RANKING place="5" resultid="1127" />
                    <RANKING place="1" resultid="1132" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11" agemax="-1" agemin="12" name="Internationale offene Wertung">
                  <RANKINGS>
                    <RANKING place="3" resultid="59" />
                    <RANKING place="7" resultid="107" />
                    <RANKING place="5" resultid="228" />
                    <RANKING place="2" resultid="934" />
                    <RANKING place="4" resultid="982" />
                    <RANKING place="6" resultid="1127" />
                    <RANKING place="1" resultid="1132" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="10" number="304" gender="M" round="FIN">
              <SWIMSTYLE stroke="SURFACE" relaycount="1" distance="1500" />
              <FEE value="650" currency="EUR" />
              <HEATS>
                <HEAT heatid="10001" number="1" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="4" agemax="13" agemin="12" name="Kategorie D" />
                <AGEGROUP agegroupid="3" agemax="15" agemin="14" name="Kategorie C">
                  <RANKINGS>
                    <RANKING place="1" resultid="122" />
                    <RANKING place="2" resultid="1323" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2" agemax="17" agemin="16" name="Kategorie B">
                  <RANKINGS>
                    <RANKING place="1" resultid="1175" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1" agemax="21" agemin="18" name="Junior:innen">
                  <RANKINGS>
                    <RANKING place="1" resultid="20" />
                    <RANKING place="3" resultid="158" />
                    <RANKING place="2" resultid="1346" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10" agemax="-1" agemin="12" name="offene Wertung">
                  <RANKINGS>
                    <RANKING place="2" resultid="20" />
                    <RANKING place="7" resultid="54" />
                    <RANKING place="6" resultid="122" />
                    <RANKING place="4" resultid="158" />
                    <RANKING place="1" resultid="930" />
                    <RANKING place="5" resultid="1175" />
                    <RANKING place="8" resultid="1323" />
                    <RANKING place="3" resultid="1346" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="11" number="5" gender="F" round="TIM">
              <SWIMSTYLE stroke="SURFACE" relaycount="4" distance="200" />
              <FEE value="1000" currency="EUR" />
              <HEATS>
                <HEAT heatid="11001" number="1" />
                <HEAT heatid="11002" number="2" />
                <HEAT heatid="11003" number="3" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="4" agemax="13" agemin="12" name="Kategorie D">
                  <RANKINGS>
                    <RANKING place="1" resultid="814" />
                    <RANKING place="2" resultid="1336" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3" agemax="15" agemin="14" name="Kategorie C">
                  <RANKINGS>
                    <RANKING place="1" resultid="249" />
                    <RANKING place="2" resultid="562" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2" agemax="17" agemin="16" name="Kategorie B">
                  <RANKINGS>
                    <RANKING place="4" resultid="358" />
                    <RANKING place="2" resultid="406" />
                    <RANKING place="3" resultid="1114" />
                    <RANKING place="1" resultid="1329" />
                    <RANKING place="5" resultid="1332" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1" agemax="21" agemin="18" name="Junior:innen">
                  <RANKINGS>
                    <RANKING place="3" resultid="502" />
                    <RANKING place="2" resultid="815" />
                    <RANKING place="1" resultid="1111" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="-1" agemin="176" easy.ak="176" calculate="TOTAL" name="Master I" />
                <AGEGROUP agegroupid="6" agemax="-1" agemin="399" easy.ak="399" calculate="TOTAL" name="Master II" />
                <AGEGROUP agegroupid="10" agemax="-1" agemin="12" name="offene Wertung">
                  <RANKINGS>
                    <RANKING place="7" resultid="133" />
                    <RANKING place="9" resultid="249" />
                    <RANKING place="11" resultid="358" />
                    <RANKING place="4" resultid="406" />
                    <RANKING place="8" resultid="502" />
                    <RANKING place="10" resultid="562" />
                    <RANKING place="2" resultid="742" />
                    <RANKING place="14" resultid="814" />
                    <RANKING place="5" resultid="815" />
                    <RANKING place="13" resultid="911" />
                    <RANKING place="1" resultid="1111" />
                    <RANKING place="6" resultid="1114" />
                    <RANKING place="3" resultid="1329" />
                    <RANKING place="12" resultid="1332" />
                    <RANKING place="15" resultid="1336" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11" agemax="-1" agemin="12" name="Internationale offene Wertung">
                  <RANKINGS>
                    <RANKING place="8" resultid="133" />
                    <RANKING place="10" resultid="249" />
                    <RANKING place="12" resultid="358" />
                    <RANKING place="5" resultid="406" />
                    <RANKING place="9" resultid="502" />
                    <RANKING place="11" resultid="562" />
                    <RANKING place="2" resultid="742" />
                    <RANKING place="15" resultid="814" />
                    <RANKING place="6" resultid="815" />
                    <RANKING place="3" resultid="907" />
                    <RANKING place="14" resultid="911" />
                    <RANKING place="1" resultid="1111" />
                    <RANKING place="7" resultid="1114" />
                    <RANKING place="4" resultid="1329" />
                    <RANKING place="13" resultid="1332" />
                    <RANKING place="16" resultid="1336" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="12" number="6" gender="M" round="TIM">
              <SWIMSTYLE stroke="SURFACE" relaycount="4" distance="200" />
              <FEE value="1000" currency="EUR" />
              <HEATS>
                <HEAT heatid="12001" number="1" />
                <HEAT heatid="12002" number="2" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="4" agemax="13" agemin="12" name="Kategorie D">
                  <RANKINGS>
                    <RANKING place="1" resultid="564" />
                    <RANKING place="2" resultid="1080" />
                    <RANKING place="3" resultid="1334" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3" agemax="15" agemin="14" name="Kategorie C">
                  <RANKINGS>
                    <RANKING place="1" resultid="90" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2" agemax="17" agemin="16" name="Kategorie B">
                  <RANKINGS>
                    <RANKING place="1" resultid="667" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1" agemax="21" agemin="18" name="Junior:innen">
                  <RANKINGS>
                    <RANKING place="3" resultid="251" />
                    <RANKING place="2" resultid="404" />
                    <RANKING place="1" resultid="1326" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="-1" agemin="176" easy.ak="176" calculate="TOTAL" name="Master I" />
                <AGEGROUP agegroupid="6" agemax="-1" agemin="399" easy.ak="399" calculate="TOTAL" name="Master II" />
                <AGEGROUP agegroupid="10" agemax="-1" agemin="12" name="offene Wertung">
                  <RANKINGS>
                    <RANKING place="7" resultid="90" />
                    <RANKING place="5" resultid="251" />
                    <RANKING place="4" resultid="404" />
                    <RANKING place="8" resultid="564" />
                    <RANKING place="6" resultid="667" />
                    <RANKING place="1" resultid="904" />
                    <RANKING place="9" resultid="1080" />
                    <RANKING place="3" resultid="1109" />
                    <RANKING place="2" resultid="1326" />
                    <RANKING place="10" resultid="1334" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
          </EVENTS>
        </SESSION>
        <SESSION number="2" date="2023-05-13" daytime="09:30" officialmeeting="08:45" warmupfrom="08:00">
          <EVENTS>
            <EVENT eventid="13" number="7" gender="F" round="PRE">
              <SWIMSTYLE stroke="IMMERSION" technique="DIVE" relaycount="1" distance="100" />
              <FEE value="650" currency="EUR" />
              <HEATS>
                <HEAT heatid="13001" number="1" />
                <HEAT heatid="13002" number="2" />
                <HEAT heatid="13003" number="3" />
                <HEAT heatid="13004" number="4" />
                <HEAT heatid="13005" number="5" />
                <HEAT heatid="13006" number="6" />
                <HEAT heatid="13007" number="7" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="4" agemax="13" agemin="12" name="Kategorie D">
                  <RANKINGS>
                    <RANKING place="9" resultid="235" />
                    <RANKING place="5" resultid="240" />
                    <RANKING place="4" resultid="361" />
                    <RANKING place="8" resultid="372" />
                    <RANKING place="5" resultid="493" />
                    <RANKING place="1" resultid="571" />
                    <RANKING place="2" resultid="726" />
                    <RANKING place="3" resultid="1074" />
                    <RANKING place="7" resultid="1387" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3" agemax="15" agemin="14" name="Kategorie C">
                  <RANKINGS>
                    <RANKING place="12" resultid="154" />
                    <RANKING place="11" resultid="223" />
                    <RANKING place="8" resultid="274" />
                    <RANKING place="10" resultid="285" />
                    <RANKING place="13" resultid="312" />
                    <RANKING place="7" resultid="377" />
                    <RANKING place="6" resultid="489" />
                    <RANKING place="5" resultid="531" />
                    <RANKING place="4" resultid="586" />
                    <RANKING place="2" resultid="1029" />
                    <RANKING place="1" resultid="1230" />
                    <RANKING place="3" resultid="1268" />
                    <RANKING place="9" resultid="1283" />
                    <RANKING place="14" resultid="1356" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2" agemax="17" agemin="16" name="Kategorie B">
                  <RANKINGS>
                    <RANKING place="5" resultid="52" />
                    <RANKING place="10" resultid="144" />
                    <RANKING place="9" resultid="382" />
                    <RANKING place="8" resultid="434" />
                    <RANKING place="2" resultid="442" />
                    <RANKING place="4" resultid="484" />
                    <RANKING place="6" resultid="625" />
                    <RANKING place="3" resultid="897" />
                    <RANKING place="7" resultid="957" />
                    <RANKING place="1" resultid="1343" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1" agemax="21" agemin="18" name="Junior:innen">
                  <RANKINGS>
                    <RANKING place="8" resultid="148" />
                    <RANKING place="1" resultid="245" />
                    <RANKING place="6" resultid="256" />
                    <RANKING place="5" resultid="294" />
                    <RANKING place="2" resultid="745" />
                    <RANKING place="3" resultid="759" />
                    <RANKING place="9" resultid="883" />
                    <RANKING place="10" resultid="1034" />
                    <RANKING place="4" resultid="1046" />
                    <RANKING place="7" resultid="1061" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="34" agemin="29" name="Master A">
                  <RANKINGS>
                    <RANKING place="1" resultid="4" />
                    <RANKING place="2" resultid="47" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6" agemax="44" agemin="35" name="Master B">
                  <RANKINGS>
                    <RANKING place="1" resultid="773" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7" agemax="54" agemin="45" name="Master C">
                  <RANKINGS>
                    <RANKING place="1" resultid="27" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8" agemax="64" agemin="55" name="Master D" />
                <AGEGROUP agegroupid="9" agemax="-1" agemin="65" name="Master E" />
                <AGEGROUP agegroupid="10" agemax="-1" agemin="12" name="offene Wertung">
                  <RANKINGS>
                    <RANKING place="20" resultid="4" />
                    <RANKING place="13" resultid="27" />
                    <RANKING place="46" resultid="47" />
                    <RANKING place="22" resultid="52" />
                    <RANKING place="8" resultid="71" />
                    <RANKING place="41" resultid="144" />
                    <RANKING place="15" resultid="148" />
                    <RANKING place="45" resultid="154" />
                    <RANKING place="44" resultid="223" />
                    <RANKING place="51" resultid="235" />
                    <RANKING place="42" resultid="240" />
                    <RANKING place="4" resultid="245" />
                    <RANKING place="12" resultid="256" />
                    <RANKING place="33" resultid="274" />
                    <RANKING place="36" resultid="285" />
                    <RANKING place="27" resultid="289" />
                    <RANKING place="11" resultid="294" />
                    <RANKING place="48" resultid="312" />
                    <RANKING place="40" resultid="361" />
                    <RANKING place="49" resultid="372" />
                    <RANKING place="30" resultid="377" />
                    <RANKING place="32" resultid="382" />
                    <RANKING place="31" resultid="434" />
                    <RANKING place="7" resultid="442" />
                    <RANKING place="19" resultid="484" />
                    <RANKING place="29" resultid="489" />
                    <RANKING place="42" resultid="493" />
                    <RANKING place="28" resultid="531" />
                    <RANKING place="24" resultid="571" />
                    <RANKING place="25" resultid="586" />
                    <RANKING place="23" resultid="625" />
                    <RANKING place="37" resultid="726" />
                    <RANKING place="5" resultid="745" />
                    <RANKING place="6" resultid="759" />
                    <RANKING place="38" resultid="773" />
                    <RANKING place="2" resultid="778" />
                    <RANKING place="17" resultid="883" />
                    <RANKING place="18" resultid="897" />
                    <RANKING place="26" resultid="957" />
                    <RANKING place="9" resultid="1029" />
                    <RANKING place="21" resultid="1034" />
                    <RANKING place="10" resultid="1046" />
                    <RANKING place="14" resultid="1061" />
                    <RANKING place="39" resultid="1074" />
                    <RANKING place="34" resultid="1156" />
                    <RANKING place="3" resultid="1230" />
                    <RANKING place="16" resultid="1268" />
                    <RANKING place="35" resultid="1283" />
                    <RANKING place="1" resultid="1343" />
                    <RANKING place="50" resultid="1356" />
                    <RANKING place="47" resultid="1387" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11" agemax="-1" agemin="12" name="Internationale Wertung">
                  <RANKINGS>
                    <RANKING place="23" resultid="4" />
                    <RANKING place="15" resultid="27" />
                    <RANKING place="17" resultid="40" />
                    <RANKING place="49" resultid="47" />
                    <RANKING place="25" resultid="52" />
                    <RANKING place="9" resultid="71" />
                    <RANKING place="44" resultid="144" />
                    <RANKING place="18" resultid="148" />
                    <RANKING place="48" resultid="154" />
                    <RANKING place="47" resultid="223" />
                    <RANKING place="55" resultid="235" />
                    <RANKING place="45" resultid="240" />
                    <RANKING place="4" resultid="245" />
                    <RANKING place="14" resultid="256" />
                    <RANKING place="36" resultid="274" />
                    <RANKING place="39" resultid="285" />
                    <RANKING place="30" resultid="289" />
                    <RANKING place="13" resultid="294" />
                    <RANKING place="52" resultid="312" />
                    <RANKING place="43" resultid="361" />
                    <RANKING place="53" resultid="372" />
                    <RANKING place="33" resultid="377" />
                    <RANKING place="35" resultid="382" />
                    <RANKING place="34" resultid="434" />
                    <RANKING place="8" resultid="442" />
                    <RANKING place="22" resultid="484" />
                    <RANKING place="32" resultid="489" />
                    <RANKING place="45" resultid="493" />
                    <RANKING place="31" resultid="531" />
                    <RANKING place="27" resultid="571" />
                    <RANKING place="28" resultid="586" />
                    <RANKING place="26" resultid="625" />
                    <RANKING place="40" resultid="726" />
                    <RANKING place="5" resultid="745" />
                    <RANKING place="6" resultid="759" />
                    <RANKING place="41" resultid="773" />
                    <RANKING place="2" resultid="778" />
                    <RANKING place="20" resultid="883" />
                    <RANKING place="21" resultid="897" />
                    <RANKING place="29" resultid="957" />
                    <RANKING place="7" resultid="961" />
                    <RANKING place="50" resultid="979" />
                    <RANKING place="11" resultid="983" />
                    <RANKING place="10" resultid="1029" />
                    <RANKING place="24" resultid="1034" />
                    <RANKING place="12" resultid="1046" />
                    <RANKING place="16" resultid="1061" />
                    <RANKING place="42" resultid="1074" />
                    <RANKING place="37" resultid="1156" />
                    <RANKING place="3" resultid="1230" />
                    <RANKING place="19" resultid="1268" />
                    <RANKING place="38" resultid="1283" />
                    <RANKING place="1" resultid="1343" />
                    <RANKING place="54" resultid="1356" />
                    <RANKING place="51" resultid="1387" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="14" number="8" gender="M" round="PRE">
              <SWIMSTYLE stroke="IMMERSION" technique="DIVE" relaycount="1" distance="100" />
              <FEE value="650" currency="EUR" />
              <HEATS>
                <HEAT heatid="14001" number="1" />
                <HEAT heatid="14002" number="2" />
                <HEAT heatid="14003" number="3" />
                <HEAT heatid="14004" number="4" />
                <HEAT heatid="14005" number="5" />
                <HEAT heatid="14006" number="6" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="4" agemax="13" agemin="12" name="Kategorie D">
                  <RANKINGS>
                    <RANKING place="1" resultid="267" />
                    <RANKING place="2" resultid="614" />
                    <RANKING place="3" resultid="673" />
                    <RANKING place="5" resultid="702" />
                    <RANKING place="6" resultid="731" />
                    <RANKING place="4" resultid="1304" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3" agemax="15" agemin="14" name="Kategorie C">
                  <RANKINGS>
                    <RANKING place="6" resultid="123" />
                    <RANKING place="4" resultid="135" />
                    <RANKING place="3" resultid="507" />
                    <RANKING place="5" resultid="523" />
                    <RANKING place="1" resultid="716" />
                    <RANKING place="2" resultid="1351" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2" agemax="17" agemin="16" name="Kategorie B">
                  <RANKINGS>
                    <RANKING place="9" resultid="99" />
                    <RANKING place="3" resultid="262" />
                    <RANKING place="1" resultid="634" />
                    <RANKING place="8" resultid="685" />
                    <RANKING place="5" resultid="721" />
                    <RANKING place="2" resultid="796" />
                    <RANKING place="6" resultid="1082" />
                    <RANKING place="4" resultid="1118" />
                    <RANKING place="7" resultid="1370" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1" agemax="21" agemin="18" name="Junior:innen">
                  <RANKINGS>
                    <RANKING place="4" resultid="21" />
                    <RANKING place="7" resultid="159" />
                    <RANKING place="5" resultid="317" />
                    <RANKING place="1" resultid="475" />
                    <RANKING place="2" resultid="690" />
                    <RANKING place="9" resultid="711" />
                    <RANKING place="8" resultid="861" />
                    <RANKING place="3" resultid="1221" />
                    <RANKING place="6" resultid="1261" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="34" agemin="29" name="Master A">
                  <RANKINGS>
                    <RANKING place="1" resultid="966" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6" agemax="44" agemin="35" name="Master B">
                  <RANKINGS>
                    <RANKING place="1" resultid="64" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7" agemax="54" agemin="45" name="Master C">
                  <RANKINGS>
                    <RANKING place="2" resultid="180" />
                    <RANKING place="3" resultid="609" />
                    <RANKING place="4" resultid="644" />
                    <RANKING place="1" resultid="783" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8" agemax="64" agemin="55" name="Master D">
                  <RANKINGS>
                    <RANKING place="1" resultid="10" />
                    <RANKING place="3" resultid="55" />
                    <RANKING place="2" resultid="199" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9" agemax="-1" agemin="65" name="Master E">
                  <RANKINGS>
                    <RANKING place="1" resultid="193" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10" agemax="-1" agemin="12" name="offene Wertung">
                  <RANKINGS>
                    <RANKING place="15" resultid="10" />
                    <RANKING place="9" resultid="21" />
                    <RANKING place="37" resultid="55" />
                    <RANKING place="14" resultid="64" />
                    <RANKING place="35" resultid="99" />
                    <RANKING place="39" resultid="123" />
                    <RANKING place="32" resultid="135" />
                    <RANKING place="18" resultid="159" />
                    <RANKING place="26" resultid="180" />
                    <RANKING place="38" resultid="193" />
                    <RANKING place="29" resultid="199" />
                    <RANKING place="19" resultid="262" />
                    <RANKING place="33" resultid="267" />
                    <RANKING place="13" resultid="317" />
                    <RANKING place="5" resultid="475" />
                    <RANKING place="30" resultid="507" />
                    <RANKING place="34" resultid="523" />
                    <RANKING place="11" resultid="557" />
                    <RANKING place="27" resultid="609" />
                    <RANKING place="36" resultid="614" />
                    <RANKING place="2" resultid="634" />
                    <RANKING place="42" resultid="644" />
                    <RANKING place="40" resultid="673" />
                    <RANKING place="31" resultid="685" />
                    <RANKING place="7" resultid="690" />
                    <RANKING place="43" resultid="702" />
                    <RANKING place="25" resultid="711" />
                    <RANKING place="10" resultid="716" />
                    <RANKING place="21" resultid="721" />
                    <RANKING place="44" resultid="731" />
                    <RANKING place="24" resultid="783" />
                    <RANKING place="3" resultid="796" />
                    <RANKING place="22" resultid="861" />
                    <RANKING place="1" resultid="946" />
                    <RANKING place="4" resultid="966" />
                    <RANKING place="23" resultid="1082" />
                    <RANKING place="20" resultid="1118" />
                    <RANKING place="12" resultid="1122" />
                    <RANKING place="8" resultid="1221" />
                    <RANKING place="17" resultid="1261" />
                    <RANKING place="41" resultid="1304" />
                    <RANKING place="16" resultid="1351" />
                    <RANKING place="6" resultid="1359" />
                    <RANKING place="28" resultid="1370" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11" agemax="-1" agemin="12" name="Internationale offene Wertung">
                  <RANKINGS>
                    <RANKING place="18" resultid="10" />
                    <RANKING place="10" resultid="21" />
                    <RANKING place="40" resultid="55" />
                    <RANKING place="17" resultid="64" />
                    <RANKING place="38" resultid="99" />
                    <RANKING place="42" resultid="123" />
                    <RANKING place="35" resultid="135" />
                    <RANKING place="21" resultid="159" />
                    <RANKING place="15" resultid="163" />
                    <RANKING place="16" resultid="167" />
                    <RANKING place="29" resultid="180" />
                    <RANKING place="41" resultid="193" />
                    <RANKING place="32" resultid="199" />
                    <RANKING place="22" resultid="262" />
                    <RANKING place="36" resultid="267" />
                    <RANKING place="14" resultid="317" />
                    <RANKING place="5" resultid="475" />
                    <RANKING place="33" resultid="507" />
                    <RANKING place="37" resultid="523" />
                    <RANKING place="12" resultid="557" />
                    <RANKING place="30" resultid="609" />
                    <RANKING place="39" resultid="614" />
                    <RANKING place="2" resultid="634" />
                    <RANKING place="45" resultid="644" />
                    <RANKING place="43" resultid="673" />
                    <RANKING place="34" resultid="685" />
                    <RANKING place="8" resultid="690" />
                    <RANKING place="46" resultid="702" />
                    <RANKING place="28" resultid="711" />
                    <RANKING place="11" resultid="716" />
                    <RANKING place="24" resultid="721" />
                    <RANKING place="47" resultid="731" />
                    <RANKING place="27" resultid="783" />
                    <RANKING place="3" resultid="796" />
                    <RANKING place="25" resultid="861" />
                    <RANKING place="1" resultid="946" />
                    <RANKING place="4" resultid="966" />
                    <RANKING place="26" resultid="1082" />
                    <RANKING place="23" resultid="1118" />
                    <RANKING place="13" resultid="1122" />
                    <RANKING place="9" resultid="1221" />
                    <RANKING place="20" resultid="1261" />
                    <RANKING place="44" resultid="1304" />
                    <RANKING place="19" resultid="1351" />
                    <RANKING place="7" resultid="1359" />
                    <RANKING place="31" resultid="1370" />
                    <RANKING place="6" resultid="1385" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="15" number="9" gender="F" round="PRE">
              <SWIMSTYLE stroke="SURFACE" relaycount="1" distance="200" />
              <FEE value="650" currency="EUR" />
              <HEATS>
                <HEAT heatid="15001" number="1" />
                <HEAT heatid="15002" number="2" />
                <HEAT heatid="15003" number="3" />
                <HEAT heatid="15004" number="4" />
                <HEAT heatid="15005" number="5" />
                <HEAT heatid="15006" number="6" />
                <HEAT heatid="15007" number="7" />
                <HEAT heatid="15008" number="8" />
                <HEAT heatid="15009" number="9" />
                <HEAT heatid="15010" number="10" />
                <HEAT heatid="15011" number="11" />
                <HEAT heatid="15012" number="12" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="4" agemax="13" agemin="12" name="Kategorie D">
                  <RANKINGS>
                    <RANKING place="11" resultid="236" />
                    <RANKING place="9" resultid="241" />
                    <RANKING place="17" resultid="304" />
                    <RANKING place="18" resultid="546" />
                    <RANKING place="1" resultid="572" />
                    <RANKING place="14" resultid="594" />
                    <RANKING place="6" resultid="669" />
                    <RANKING place="5" resultid="727" />
                    <RANKING place="16" resultid="788" />
                    <RANKING place="8" resultid="792" />
                    <RANKING place="2" resultid="823" />
                    <RANKING place="13" resultid="833" />
                    <RANKING place="3" resultid="872" />
                    <RANKING place="4" resultid="878" />
                    <RANKING place="10" resultid="944" />
                    <RANKING place="12" resultid="1054" />
                    <RANKING place="15" resultid="1075" />
                    <RANKING place="19" resultid="1288" />
                    <RANKING place="7" resultid="1295" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3" agemax="15" agemin="14" name="Kategorie C">
                  <RANKINGS>
                    <RANKING place="16" resultid="155" />
                    <RANKING place="20" resultid="224" />
                    <RANKING place="9" resultid="275" />
                    <RANKING place="7" resultid="281" />
                    <RANKING place="17" resultid="313" />
                    <RANKING place="13" resultid="412" />
                    <RANKING place="10" resultid="438" />
                    <RANKING place="2" resultid="465" />
                    <RANKING place="6" resultid="587" />
                    <RANKING place="21" resultid="598" />
                    <RANKING place="14" resultid="640" />
                    <RANKING place="12" resultid="842" />
                    <RANKING place="4" resultid="953" />
                    <RANKING place="5" resultid="1206" />
                    <RANKING place="3" resultid="1211" />
                    <RANKING place="1" resultid="1231" />
                    <RANKING place="23" resultid="1236" />
                    <RANKING place="8" resultid="1269" />
                    <RANKING place="18" resultid="1277" />
                    <RANKING place="11" resultid="1284" />
                    <RANKING place="19" resultid="1315" />
                    <RANKING place="22" resultid="1357" />
                    <RANKING place="15" resultid="1364" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2" agemax="17" agemin="16" name="Kategorie B">
                  <RANKINGS>
                    <RANKING place="6" resultid="229" />
                    <RANKING place="1" resultid="425" />
                    <RANKING place="4" resultid="443" />
                    <RANKING place="14" resultid="518" />
                    <RANKING place="12" resultid="626" />
                    <RANKING place="11" resultid="898" />
                    <RANKING place="2" resultid="935" />
                    <RANKING place="8" resultid="1097" />
                    <RANKING place="9" resultid="1101" />
                    <RANKING place="5" resultid="1139" />
                    <RANKING place="10" resultid="1148" />
                    <RANKING place="15" resultid="1152" />
                    <RANKING place="3" resultid="1165" />
                    <RANKING place="13" resultid="1225" />
                    <RANKING place="7" resultid="1309" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1" agemax="21" agemin="18" name="Junior:innen">
                  <RANKINGS>
                    <RANKING place="7" resultid="76" />
                    <RANKING place="12" resultid="108" />
                    <RANKING place="4" resultid="246" />
                    <RANKING place="11" resultid="257" />
                    <RANKING place="9" resultid="295" />
                    <RANKING place="8" resultid="535" />
                    <RANKING place="6" resultid="767" />
                    <RANKING place="5" resultid="866" />
                    <RANKING place="3" resultid="975" />
                    <RANKING place="10" resultid="1128" />
                    <RANKING place="1" resultid="1133" />
                    <RANKING place="2" resultid="1144" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="34" agemin="29" name="Master A">
                  <RANKINGS>
                    <RANKING place="1" resultid="5" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6" agemax="44" agemin="35" name="Master B">
                  <RANKINGS>
                    <RANKING place="1" resultid="648" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7" agemax="54" agemin="45" name="Master C">
                  <RANKINGS>
                    <RANKING place="1" resultid="837" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8" agemax="64" agemin="55" name="Master D">
                  <RANKINGS>
                    <RANKING place="1" resultid="658" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9" agemax="-1" agemin="65" name="Master E" />
                <AGEGROUP agegroupid="10" agemax="-1" agemin="12" name="offene Wertung">
                  <RANKINGS>
                    <RANKING place="30" resultid="5" />
                    <RANKING place="16" resultid="60" />
                    <RANKING place="13" resultid="76" />
                    <RANKING place="10" resultid="83" />
                    <RANKING place="33" resultid="108" />
                    <RANKING place="35" resultid="117" />
                    <RANKING place="34" resultid="141" />
                    <RANKING place="58" resultid="155" />
                    <RANKING place="67" resultid="224" />
                    <RANKING place="22" resultid="229" />
                    <RANKING place="71" resultid="236" />
                    <RANKING place="65" resultid="241" />
                    <RANKING place="5" resultid="246" />
                    <RANKING place="27" resultid="257" />
                    <RANKING place="44" resultid="275" />
                    <RANKING place="42" resultid="281" />
                    <RANKING place="50" resultid="290" />
                    <RANKING place="19" resultid="295" />
                    <RANKING place="78" resultid="304" />
                    <RANKING place="59" resultid="313" />
                    <RANKING place="52" resultid="412" />
                    <RANKING place="6" resultid="425" />
                    <RANKING place="45" resultid="438" />
                    <RANKING place="15" resultid="443" />
                    <RANKING place="18" resultid="465" />
                    <RANKING place="48" resultid="518" />
                    <RANKING place="17" resultid="535" />
                    <RANKING place="79" resultid="546" />
                    <RANKING place="32" resultid="572" />
                    <RANKING place="38" resultid="587" />
                    <RANKING place="75" resultid="594" />
                    <RANKING place="68" resultid="598" />
                    <RANKING place="40" resultid="626" />
                    <RANKING place="54" resultid="640" />
                    <RANKING place="53" resultid="648" />
                    <RANKING place="81" resultid="658" />
                    <RANKING place="62" resultid="669" />
                    <RANKING place="60" resultid="727" />
                    <RANKING place="12" resultid="767" />
                    <RANKING place="2" resultid="779" />
                    <RANKING place="77" resultid="788" />
                    <RANKING place="64" resultid="792" />
                    <RANKING place="39" resultid="823" />
                    <RANKING place="74" resultid="833" />
                    <RANKING place="47" resultid="837" />
                    <RANKING place="51" resultid="842" />
                    <RANKING place="11" resultid="866" />
                    <RANKING place="41" resultid="872" />
                    <RANKING place="56" resultid="878" />
                    <RANKING place="37" resultid="898" />
                    <RANKING place="28" resultid="928" />
                    <RANKING place="7" resultid="935" />
                    <RANKING place="70" resultid="944" />
                    <RANKING place="25" resultid="953" />
                    <RANKING place="4" resultid="975" />
                    <RANKING place="73" resultid="1054" />
                    <RANKING place="76" resultid="1075" />
                    <RANKING place="26" resultid="1097" />
                    <RANKING place="29" resultid="1101" />
                    <RANKING place="21" resultid="1128" />
                    <RANKING place="1" resultid="1133" />
                    <RANKING place="20" resultid="1139" />
                    <RANKING place="3" resultid="1144" />
                    <RANKING place="31" resultid="1148" />
                    <RANKING place="55" resultid="1152" />
                    <RANKING place="14" resultid="1165" />
                    <RANKING place="36" resultid="1206" />
                    <RANKING place="23" resultid="1211" />
                    <RANKING place="46" resultid="1225" />
                    <RANKING place="8" resultid="1231" />
                    <RANKING place="72" resultid="1236" />
                    <RANKING place="43" resultid="1269" />
                    <RANKING place="61" resultid="1277" />
                    <RANKING place="49" resultid="1284" />
                    <RANKING place="80" resultid="1288" />
                    <RANKING place="63" resultid="1295" />
                    <RANKING place="9" resultid="1301" />
                    <RANKING place="24" resultid="1309" />
                    <RANKING place="66" resultid="1315" />
                    <RANKING place="69" resultid="1357" />
                    <RANKING place="57" resultid="1364" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11" agemax="-1" agemin="12" name="Internationale offene Wertung">
                  <RANKINGS>
                    <RANKING place="32" resultid="5" />
                    <RANKING place="18" resultid="60" />
                    <RANKING place="14" resultid="76" />
                    <RANKING place="11" resultid="83" />
                    <RANKING place="36" resultid="108" />
                    <RANKING place="38" resultid="117" />
                    <RANKING place="37" resultid="141" />
                    <RANKING place="63" resultid="155" />
                    <RANKING place="71" resultid="214" />
                    <RANKING place="73" resultid="224" />
                    <RANKING place="24" resultid="229" />
                    <RANKING place="77" resultid="236" />
                    <RANKING place="70" resultid="241" />
                    <RANKING place="5" resultid="246" />
                    <RANKING place="29" resultid="257" />
                    <RANKING place="47" resultid="275" />
                    <RANKING place="45" resultid="281" />
                    <RANKING place="54" resultid="290" />
                    <RANKING place="21" resultid="295" />
                    <RANKING place="84" resultid="304" />
                    <RANKING place="64" resultid="313" />
                    <RANKING place="56" resultid="412" />
                    <RANKING place="7" resultid="425" />
                    <RANKING place="48" resultid="438" />
                    <RANKING place="17" resultid="443" />
                    <RANKING place="60" resultid="460" />
                    <RANKING place="20" resultid="465" />
                    <RANKING place="52" resultid="518" />
                    <RANKING place="19" resultid="535" />
                    <RANKING place="85" resultid="546" />
                    <RANKING place="35" resultid="572" />
                    <RANKING place="34" resultid="576" />
                    <RANKING place="41" resultid="587" />
                    <RANKING place="81" resultid="594" />
                    <RANKING place="74" resultid="598" />
                    <RANKING place="43" resultid="626" />
                    <RANKING place="58" resultid="640" />
                    <RANKING place="57" resultid="648" />
                    <RANKING place="87" resultid="658" />
                    <RANKING place="67" resultid="669" />
                    <RANKING place="49" resultid="708" />
                    <RANKING place="65" resultid="727" />
                    <RANKING place="13" resultid="767" />
                    <RANKING place="2" resultid="779" />
                    <RANKING place="83" resultid="788" />
                    <RANKING place="69" resultid="792" />
                    <RANKING place="42" resultid="823" />
                    <RANKING place="80" resultid="833" />
                    <RANKING place="51" resultid="837" />
                    <RANKING place="55" resultid="842" />
                    <RANKING place="12" resultid="866" />
                    <RANKING place="44" resultid="872" />
                    <RANKING place="61" resultid="878" />
                    <RANKING place="40" resultid="898" />
                    <RANKING place="30" resultid="928" />
                    <RANKING place="8" resultid="935" />
                    <RANKING place="76" resultid="944" />
                    <RANKING place="27" resultid="953" />
                    <RANKING place="6" resultid="962" />
                    <RANKING place="4" resultid="975" />
                    <RANKING place="79" resultid="1054" />
                    <RANKING place="82" resultid="1075" />
                    <RANKING place="28" resultid="1097" />
                    <RANKING place="31" resultid="1101" />
                    <RANKING place="23" resultid="1128" />
                    <RANKING place="1" resultid="1133" />
                    <RANKING place="22" resultid="1139" />
                    <RANKING place="3" resultid="1144" />
                    <RANKING place="33" resultid="1148" />
                    <RANKING place="59" resultid="1152" />
                    <RANKING place="16" resultid="1159" />
                    <RANKING place="15" resultid="1165" />
                    <RANKING place="39" resultid="1206" />
                    <RANKING place="25" resultid="1211" />
                    <RANKING place="50" resultid="1225" />
                    <RANKING place="9" resultid="1231" />
                    <RANKING place="78" resultid="1236" />
                    <RANKING place="46" resultid="1269" />
                    <RANKING place="66" resultid="1277" />
                    <RANKING place="53" resultid="1284" />
                    <RANKING place="86" resultid="1288" />
                    <RANKING place="68" resultid="1295" />
                    <RANKING place="10" resultid="1301" />
                    <RANKING place="26" resultid="1309" />
                    <RANKING place="72" resultid="1315" />
                    <RANKING place="75" resultid="1357" />
                    <RANKING place="62" resultid="1364" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="16" number="10" gender="M" round="PRE">
              <SWIMSTYLE stroke="SURFACE" relaycount="1" distance="200" />
              <FEE value="650" currency="EUR" />
              <HEATS>
                <HEAT heatid="16001" number="1" />
                <HEAT heatid="16002" number="2" />
                <HEAT heatid="16003" number="3" />
                <HEAT heatid="16004" number="4" />
                <HEAT heatid="16005" number="5" />
                <HEAT heatid="16006" number="6" />
                <HEAT heatid="16007" number="7" />
                <HEAT heatid="16008" number="8" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="4" agemax="13" agemin="12" name="Kategorie D">
                  <RANKINGS>
                    <RANKING place="8" resultid="94" />
                    <RANKING place="2" resultid="268" />
                    <RANKING place="11" resultid="591" />
                    <RANKING place="1" resultid="615" />
                    <RANKING place="7" resultid="621" />
                    <RANKING place="10" resultid="631" />
                    <RANKING place="6" resultid="674" />
                    <RANKING place="3" resultid="703" />
                    <RANKING place="9" resultid="732" />
                    <RANKING place="5" resultid="1090" />
                    <RANKING place="12" resultid="1188" />
                    <RANKING place="13" resultid="1299" />
                    <RANKING place="4" resultid="1305" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3" agemax="15" agemin="14" name="Kategorie C">
                  <RANKINGS>
                    <RANKING place="16" resultid="113" />
                    <RANKING place="9" resultid="124" />
                    <RANKING place="15" resultid="128" />
                    <RANKING place="8" resultid="136" />
                    <RANKING place="11" resultid="398" />
                    <RANKING place="1" resultid="416" />
                    <RANKING place="5" resultid="449" />
                    <RANKING place="12" resultid="508" />
                    <RANKING place="3" resultid="528" />
                    <RANKING place="10" resultid="601" />
                    <RANKING place="14" resultid="605" />
                    <RANKING place="17" resultid="849" />
                    <RANKING place="4" resultid="916" />
                    <RANKING place="7" resultid="1085" />
                    <RANKING place="6" resultid="1197" />
                    <RANKING place="13" resultid="1217" />
                    <RANKING place="2" resultid="1352" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2" agemax="17" agemin="16" name="Kategorie B">
                  <RANKINGS>
                    <RANKING place="7" resultid="100" />
                    <RANKING place="4" resultid="263" />
                    <RANKING place="1" resultid="635" />
                    <RANKING place="2" resultid="797" />
                    <RANKING place="3" resultid="923" />
                    <RANKING place="6" resultid="1119" />
                    <RANKING place="5" resultid="1176" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1" agemax="21" agemin="18" name="Junior:innen">
                  <RANKINGS>
                    <RANKING place="5" resultid="299" />
                    <RANKING place="2" resultid="387" />
                    <RANKING place="3" resultid="691" />
                    <RANKING place="4" resultid="1202" />
                    <RANKING place="1" resultid="1263" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="34" agemin="29" name="Master A">
                  <RANKINGS>
                    <RANKING place="1" resultid="967" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6" agemax="44" agemin="35" name="Master B">
                  <RANKINGS>
                    <RANKING place="2" resultid="33" />
                    <RANKING place="1" resultid="65" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7" agemax="54" agemin="45" name="Master C">
                  <RANKINGS>
                    <RANKING place="2" resultid="181" />
                    <RANKING place="3" resultid="540" />
                    <RANKING place="1" resultid="1009" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8" agemax="64" agemin="55" name="Master D">
                  <RANKINGS>
                    <RANKING place="1" resultid="11" />
                    <RANKING place="2" resultid="200" />
                    <RANKING place="4" resultid="737" />
                    <RANKING place="3" resultid="828" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9" agemax="-1" agemin="65" name="Master E">
                  <RANKINGS>
                    <RANKING place="1" resultid="752" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10" agemax="-1" agemin="12" name="offene Wertung">
                  <RANKINGS>
                    <RANKING place="25" resultid="11" />
                    <RANKING place="33" resultid="33" />
                    <RANKING place="23" resultid="65" />
                    <RANKING place="51" resultid="94" />
                    <RANKING place="29" resultid="100" />
                    <RANKING place="45" resultid="113" />
                    <RANKING place="31" resultid="124" />
                    <RANKING place="44" resultid="128" />
                    <RANKING place="30" resultid="136" />
                    <RANKING place="34" resultid="181" />
                    <RANKING place="39" resultid="200" />
                    <RANKING place="19" resultid="263" />
                    <RANKING place="40" resultid="268" />
                    <RANKING place="27" resultid="299" />
                    <RANKING place="8" resultid="387" />
                    <RANKING place="35" resultid="398" />
                    <RANKING place="13" resultid="416" />
                    <RANKING place="24" resultid="449" />
                    <RANKING place="37" resultid="508" />
                    <RANKING place="16" resultid="528" />
                    <RANKING place="41" resultid="540" />
                    <RANKING place="56" resultid="591" />
                    <RANKING place="32" resultid="601" />
                    <RANKING place="43" resultid="605" />
                    <RANKING place="35" resultid="615" />
                    <RANKING place="50" resultid="621" />
                    <RANKING place="54" resultid="631" />
                    <RANKING place="4" resultid="635" />
                    <RANKING place="49" resultid="674" />
                    <RANKING place="11" resultid="691" />
                    <RANKING place="42" resultid="703" />
                    <RANKING place="53" resultid="732" />
                    <RANKING place="55" resultid="737" />
                    <RANKING place="59" resultid="752" />
                    <RANKING place="5" resultid="797" />
                    <RANKING place="52" resultid="828" />
                    <RANKING place="46" resultid="849" />
                    <RANKING place="15" resultid="888" />
                    <RANKING place="17" resultid="916" />
                    <RANKING place="9" resultid="923" />
                    <RANKING place="3" resultid="931" />
                    <RANKING place="7" resultid="940" />
                    <RANKING place="2" resultid="947" />
                    <RANKING place="1" resultid="967" />
                    <RANKING place="20" resultid="1009" />
                    <RANKING place="28" resultid="1085" />
                    <RANKING place="48" resultid="1090" />
                    <RANKING place="22" resultid="1119" />
                    <RANKING place="12" resultid="1123" />
                    <RANKING place="21" resultid="1176" />
                    <RANKING place="57" resultid="1188" />
                    <RANKING place="26" resultid="1197" />
                    <RANKING place="18" resultid="1202" />
                    <RANKING place="38" resultid="1217" />
                    <RANKING place="6" resultid="1263" />
                    <RANKING place="58" resultid="1299" />
                    <RANKING place="47" resultid="1305" />
                    <RANKING place="14" resultid="1352" />
                    <RANKING place="10" resultid="1360" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="17" number="11" gender="F" round="TIM">
              <SWIMSTYLE stroke="SURFACE" relaycount="1" distance="800" />
              <FEE value="650" currency="EUR" />
              <HEATS>
                <HEAT heatid="17001" number="1" />
                <HEAT heatid="17002" number="2" />
                <HEAT heatid="17003" number="3" />
                <HEAT heatid="17004" number="4" />
                <HEAT heatid="17005" number="5" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="4" agemax="13" agemin="12" name="Kategorie D">
                  <RANKINGS>
                    <RANKING place="3" resultid="362" />
                    <RANKING place="7" resultid="373" />
                    <RANKING place="1" resultid="421" />
                    <RANKING place="8" resultid="547" />
                    <RANKING place="5" resultid="824" />
                    <RANKING place="2" resultid="873" />
                    <RANKING place="4" resultid="879" />
                    <RANKING place="6" resultid="1296" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3" agemax="15" agemin="14" name="Kategorie C">
                  <RANKINGS>
                    <RANKING place="1" resultid="378" />
                    <RANKING place="2" resultid="641" />
                    <RANKING place="4" resultid="843" />
                    <RANKING place="3" resultid="1365" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2" agemax="17" agemin="16" name="Kategorie B">
                  <RANKINGS>
                    <RANKING place="2" resultid="53" />
                    <RANKING place="5" resultid="230" />
                    <RANKING place="7" resultid="383" />
                    <RANKING place="4" resultid="1102" />
                    <RANKING place="3" resultid="1140" />
                    <RANKING place="1" resultid="1166" />
                    <RANKING place="8" resultid="1192" />
                    <RANKING place="6" resultid="1254" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1" agemax="21" agemin="18" name="Junior:innen">
                  <RANKINGS>
                    <RANKING place="1" resultid="109" />
                    <RANKING place="2" resultid="149" />
                    <RANKING place="3" resultid="1062" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="34" agemin="29" name="Master A">
                  <RANKINGS>
                    <RANKING place="1" resultid="6" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6" agemax="44" agemin="35" name="Master B">
                  <RANKINGS>
                    <RANKING place="1" resultid="649" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7" agemax="54" agemin="45" name="Master C">
                  <RANKINGS>
                    <RANKING place="1" resultid="28" />
                    <RANKING place="2" resultid="838" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8" agemax="64" agemin="55" name="Master D" />
                <AGEGROUP agegroupid="9" agemax="-1" agemin="65" name="Master E" />
                <AGEGROUP agegroupid="10" agemax="-1" agemin="12" name="offene Wertung">
                  <RANKINGS>
                    <RANKING place="5" resultid="6" />
                    <RANKING place="13" resultid="28" />
                    <RANKING place="2" resultid="53" />
                    <RANKING place="7" resultid="109" />
                    <RANKING place="10" resultid="118" />
                    <RANKING place="11" resultid="142" />
                    <RANKING place="9" resultid="149" />
                    <RANKING place="6" resultid="230" />
                    <RANKING place="21" resultid="362" />
                    <RANKING place="28" resultid="373" />
                    <RANKING place="15" resultid="378" />
                    <RANKING place="12" resultid="383" />
                    <RANKING place="16" resultid="421" />
                    <RANKING place="29" resultid="547" />
                    <RANKING place="18" resultid="641" />
                    <RANKING place="27" resultid="649" />
                    <RANKING place="25" resultid="824" />
                    <RANKING place="23" resultid="838" />
                    <RANKING place="24" resultid="843" />
                    <RANKING place="19" resultid="873" />
                    <RANKING place="22" resultid="879" />
                    <RANKING place="17" resultid="1062" />
                    <RANKING place="4" resultid="1102" />
                    <RANKING place="3" resultid="1140" />
                    <RANKING place="1" resultid="1166" />
                    <RANKING place="14" resultid="1192" />
                    <RANKING place="8" resultid="1254" />
                    <RANKING place="26" resultid="1296" />
                    <RANKING place="20" resultid="1365" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11" agemax="-1" agemin="12" name="Internationale Wertung">
                  <RANKINGS>
                    <RANKING place="6" resultid="6" />
                    <RANKING place="16" resultid="28" />
                    <RANKING place="7" resultid="41" />
                    <RANKING place="3" resultid="53" />
                    <RANKING place="9" resultid="109" />
                    <RANKING place="13" resultid="118" />
                    <RANKING place="14" resultid="142" />
                    <RANKING place="11" resultid="149" />
                    <RANKING place="8" resultid="230" />
                    <RANKING place="24" resultid="362" />
                    <RANKING place="31" resultid="373" />
                    <RANKING place="18" resultid="378" />
                    <RANKING place="15" resultid="383" />
                    <RANKING place="19" resultid="421" />
                    <RANKING place="32" resultid="547" />
                    <RANKING place="12" resultid="577" />
                    <RANKING place="21" resultid="641" />
                    <RANKING place="30" resultid="649" />
                    <RANKING place="28" resultid="824" />
                    <RANKING place="26" resultid="838" />
                    <RANKING place="27" resultid="843" />
                    <RANKING place="22" resultid="873" />
                    <RANKING place="25" resultid="879" />
                    <RANKING place="1" resultid="984" />
                    <RANKING place="20" resultid="1062" />
                    <RANKING place="5" resultid="1102" />
                    <RANKING place="4" resultid="1140" />
                    <RANKING place="2" resultid="1166" />
                    <RANKING place="17" resultid="1192" />
                    <RANKING place="10" resultid="1254" />
                    <RANKING place="29" resultid="1296" />
                    <RANKING place="23" resultid="1365" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="18" number="12" gender="M" round="TIM">
              <SWIMSTYLE stroke="SURFACE" relaycount="1" distance="800" />
              <FEE value="650" currency="EUR" />
              <HEATS>
                <HEAT heatid="18001" number="1" />
                <HEAT heatid="18002" number="2" />
                <HEAT heatid="18003" number="3" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="4" agemax="13" agemin="12" name="Kategorie D">
                  <RANKINGS>
                    <RANKING place="1" resultid="95" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3" agemax="15" agemin="14" name="Kategorie C">
                  <RANKINGS>
                    <RANKING place="1" resultid="125" />
                    <RANKING place="5" resultid="129" />
                    <RANKING place="4" resultid="399" />
                    <RANKING place="6" resultid="606" />
                    <RANKING place="2" resultid="1086" />
                    <RANKING place="7" resultid="1291" />
                    <RANKING place="3" resultid="1324" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2" agemax="17" agemin="16" name="Kategorie B">
                  <RANKINGS>
                    <RANKING place="1" resultid="101" />
                    <RANKING place="2" resultid="1371" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1" agemax="21" agemin="18" name="Junior:innen">
                  <RANKINGS>
                    <RANKING place="1" resultid="300" />
                    <RANKING place="2" resultid="308" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="34" agemin="29" name="Master A" />
                <AGEGROUP agegroupid="6" agemax="44" agemin="35" name="Master B">
                  <RANKINGS>
                    <RANKING place="2" resultid="34" />
                    <RANKING place="1" resultid="66" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7" agemax="54" agemin="45" name="Master C">
                  <RANKINGS>
                    <RANKING place="1" resultid="801" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8" agemax="64" agemin="55" name="Master D">
                  <RANKINGS>
                    <RANKING place="1" resultid="12" />
                    <RANKING place="2" resultid="56" />
                    <RANKING place="3" resultid="201" />
                    <RANKING place="4" resultid="738" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9" agemax="-1" agemin="65" name="Master E">
                  <RANKINGS>
                    <RANKING place="2" resultid="753" />
                    <RANKING place="1" resultid="1320" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10" agemax="-1" agemin="12" name="offene Wertung">
                  <RANKINGS>
                    <RANKING place="1" resultid="12" />
                    <RANKING place="10" resultid="34" />
                    <RANKING place="9" resultid="56" />
                    <RANKING place="3" resultid="66" />
                    <RANKING place="15" resultid="95" />
                    <RANKING place="6" resultid="101" />
                    <RANKING place="5" resultid="125" />
                    <RANKING place="14" resultid="129" />
                    <RANKING place="13" resultid="201" />
                    <RANKING place="2" resultid="300" />
                    <RANKING place="4" resultid="308" />
                    <RANKING place="12" resultid="399" />
                    <RANKING place="16" resultid="606" />
                    <RANKING place="19" resultid="738" />
                    <RANKING place="21" resultid="753" />
                    <RANKING place="17" resultid="801" />
                    <RANKING place="7" resultid="1086" />
                    <RANKING place="18" resultid="1291" />
                    <RANKING place="20" resultid="1320" />
                    <RANKING place="8" resultid="1324" />
                    <RANKING place="11" resultid="1371" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11" agemax="-1" agemin="12" name="Internationale offene Wertung">
                  <RANKINGS>
                    <RANKING place="1" resultid="12" />
                    <RANKING place="10" resultid="34" />
                    <RANKING place="9" resultid="56" />
                    <RANKING place="3" resultid="66" />
                    <RANKING place="15" resultid="95" />
                    <RANKING place="6" resultid="101" />
                    <RANKING place="5" resultid="125" />
                    <RANKING place="14" resultid="129" />
                    <RANKING place="13" resultid="201" />
                    <RANKING place="2" resultid="300" />
                    <RANKING place="4" resultid="308" />
                    <RANKING place="12" resultid="399" />
                    <RANKING place="16" resultid="606" />
                    <RANKING place="19" resultid="738" />
                    <RANKING place="21" resultid="753" />
                    <RANKING place="17" resultid="801" />
                    <RANKING place="7" resultid="1086" />
                    <RANKING place="18" resultid="1291" />
                    <RANKING place="20" resultid="1320" />
                    <RANKING place="8" resultid="1324" />
                    <RANKING place="11" resultid="1371" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="19" number="13" gender="F" round="TIM">
              <SWIMSTYLE stroke="IMMERSION" technique="DIVE" relaycount="1" distance="400" />
              <FEE value="650" currency="EUR" />
              <HEATS>
                <HEAT heatid="19001" number="1" />
                <HEAT heatid="19002" number="2" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="4" agemax="13" agemin="12" name="Kategorie D" />
                <AGEGROUP agegroupid="3" agemax="15" agemin="14" name="Kategorie C">
                  <RANKINGS>
                    <RANKING place="1" resultid="276" />
                    <RANKING place="2" resultid="532" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2" agemax="17" agemin="16" name="Kategorie B">
                  <RANKINGS>
                    <RANKING place="3" resultid="145" />
                    <RANKING place="1" resultid="485" />
                    <RANKING place="2" resultid="899" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1" agemax="21" agemin="18" name="Junior:innen">
                  <RANKINGS>
                    <RANKING place="3" resultid="150" />
                    <RANKING place="4" resultid="258" />
                    <RANKING place="1" resultid="760" />
                    <RANKING place="2" resultid="1047" />
                    <RANKING place="5" resultid="1063" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="34" agemin="29" name="Master A">
                  <RANKINGS>
                    <RANKING place="1" resultid="1380" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6" agemax="44" agemin="35" name="Master B">
                  <RANKINGS>
                    <RANKING place="1" resultid="774" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7" agemax="54" agemin="45" name="Master C">
                  <RANKINGS>
                    <RANKING place="1" resultid="29" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8" agemax="64" agemin="55" name="Master D" />
                <AGEGROUP agegroupid="9" agemax="-1" agemin="65" name="Master E" />
                <AGEGROUP agegroupid="10" agemax="-1" agemin="12" name="offene Wertung">
                  <RANKINGS>
                    <RANKING place="2" resultid="29" />
                    <RANKING place="3" resultid="84" />
                    <RANKING place="13" resultid="145" />
                    <RANKING place="5" resultid="150" />
                    <RANKING place="6" resultid="258" />
                    <RANKING place="9" resultid="276" />
                    <RANKING place="8" resultid="485" />
                    <RANKING place="10" resultid="532" />
                    <RANKING place="1" resultid="760" />
                    <RANKING place="11" resultid="774" />
                    <RANKING place="12" resultid="899" />
                    <RANKING place="4" resultid="1047" />
                    <RANKING place="7" resultid="1063" />
                    <RANKING place="14" resultid="1380" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11" agemax="-1" agemin="12" name="Internationale Wertung">
                  <RANKINGS>
                    <RANKING place="2" resultid="29" />
                    <RANKING place="3" resultid="84" />
                    <RANKING place="13" resultid="145" />
                    <RANKING place="5" resultid="150" />
                    <RANKING place="6" resultid="258" />
                    <RANKING place="9" resultid="276" />
                    <RANKING place="8" resultid="485" />
                    <RANKING place="10" resultid="532" />
                    <RANKING place="1" resultid="760" />
                    <RANKING place="11" resultid="774" />
                    <RANKING place="12" resultid="899" />
                    <RANKING place="4" resultid="1047" />
                    <RANKING place="7" resultid="1063" />
                    <RANKING place="14" resultid="1380" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="20" number="14" gender="M" round="TIM">
              <SWIMSTYLE stroke="IMMERSION" technique="DIVE" relaycount="1" distance="400" />
              <FEE value="650" currency="EUR" />
              <HEATS>
                <HEAT heatid="20001" number="1" />
                <HEAT heatid="20002" number="2" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="4" agemax="13" agemin="12" name="Kategorie D">
                  <RANKINGS>
                    <RANKING place="1" resultid="269" />
                    <RANKING place="2" resultid="616" />
                    <RANKING place="3" resultid="675" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3" agemax="15" agemin="14" name="Kategorie C">
                  <RANKINGS>
                    <RANKING place="2" resultid="137" />
                    <RANKING place="1" resultid="524" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2" agemax="17" agemin="16" name="Kategorie B">
                  <RANKINGS>
                    <RANKING place="1" resultid="1372" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1" agemax="21" agemin="18" name="Junior:innen">
                  <RANKINGS>
                    <RANKING place="1" resultid="1348" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="34" agemin="29" name="Master A" />
                <AGEGROUP agegroupid="6" agemax="44" agemin="35" name="Master B" />
                <AGEGROUP agegroupid="7" agemax="54" agemin="45" name="Master C">
                  <RANKINGS>
                    <RANKING place="2" resultid="182" />
                    <RANKING place="1" resultid="610" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8" agemax="64" agemin="55" name="Master D">
                  <RANKINGS>
                    <RANKING place="1" resultid="13" />
                    <RANKING place="2" resultid="202" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9" agemax="-1" agemin="65" name="Master E">
                  <RANKINGS>
                    <RANKING place="1" resultid="194" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10" agemax="-1" agemin="12" name="offene Wertung">
                  <RANKINGS>
                    <RANKING place="2" resultid="13" />
                    <RANKING place="9" resultid="137" />
                    <RANKING place="6" resultid="182" />
                    <RANKING place="10" resultid="194" />
                    <RANKING place="4" resultid="202" />
                    <RANKING place="8" resultid="269" />
                    <RANKING place="7" resultid="524" />
                    <RANKING place="3" resultid="610" />
                    <RANKING place="11" resultid="616" />
                    <RANKING place="12" resultid="675" />
                    <RANKING place="1" resultid="1348" />
                    <RANKING place="5" resultid="1372" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11" agemax="-1" agemin="12" name="Internationale offene Wertung">
                  <RANKINGS>
                    <RANKING place="2" resultid="13" />
                    <RANKING place="9" resultid="137" />
                    <RANKING place="6" resultid="182" />
                    <RANKING place="10" resultid="194" />
                    <RANKING place="4" resultid="202" />
                    <RANKING place="8" resultid="269" />
                    <RANKING place="7" resultid="524" />
                    <RANKING place="3" resultid="610" />
                    <RANKING place="11" resultid="616" />
                    <RANKING place="12" resultid="675" />
                    <RANKING place="1" resultid="1348" />
                    <RANKING place="5" resultid="1372" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
          </EVENTS>
        </SESSION>
        <SESSION number="3" date="2023-05-13" daytime="16:05" officialmeeting="15:30" warmupfrom="15:00">
          <EVENTS>
            <EVENT eventid="21" number="107" gender="F" round="FIN">
              <SWIMSTYLE stroke="IMMERSION" technique="DIVE" relaycount="1" distance="100" />
              <HEATS>
                <HEAT heatid="21000" number="0" />
                <HEAT heatid="21001" number="1" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="10" agemax="-1" agemin="12" name="offene Wertung">
                  <RANKINGS>
                    <RANKING place="2" resultid="1493" />
                    <RANKING place="1" resultid="1494" />
                    <RANKING place="5" resultid="1495" />
                    <RANKING place="3" resultid="1496" />
                    <RANKING place="4" resultid="1497" />
                    <RANKING place="6" resultid="1499" />
                    <RANKING place="7" resultid="1500" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11" agemax="-1" agemin="12" name="Internationale offene Wertung">
                  <RANKINGS>
                    <RANKING place="2" resultid="1493" />
                    <RANKING place="1" resultid="1494" />
                    <RANKING place="5" resultid="1495" />
                    <RANKING place="3" resultid="1496" />
                    <RANKING place="4" resultid="1497" />
                    <RANKING place="6" resultid="1498" />
                    <RANKING place="7" resultid="1499" />
                    <RANKING place="8" resultid="1500" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="22" number="108" gender="M" round="FIN">
              <SWIMSTYLE stroke="IMMERSION" technique="DIVE" relaycount="1" distance="100" />
              <HEATS>
                <HEAT heatid="22000" number="0" />
                <HEAT heatid="22001" number="1" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="10" agemax="-1" agemin="12" name="offene Wertung">
                  <RANKINGS>
                    <RANKING place="1" resultid="1504" />
                    <RANKING place="4" resultid="1505" />
                    <RANKING place="3" resultid="1506" />
                    <RANKING place="2" resultid="1507" />
                    <RANKING place="6" resultid="1508" />
                    <RANKING place="5" resultid="1509" />
                    <RANKING place="7" resultid="1510" />
                    <RANKING place="8" resultid="1511" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11" agemax="-1" agemin="12" name="Internationale offene Wertung">
                  <RANKINGS>
                    <RANKING place="1" resultid="1504" />
                    <RANKING place="4" resultid="1505" />
                    <RANKING place="3" resultid="1506" />
                    <RANKING place="2" resultid="1507" />
                    <RANKING place="6" resultid="1508" />
                    <RANKING place="5" resultid="1509" />
                    <RANKING place="7" resultid="1510" />
                    <RANKING place="8" resultid="1511" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="23" number="109" gender="F" round="FIN">
              <SWIMSTYLE stroke="SURFACE" relaycount="1" distance="200" />
              <HEATS>
                <HEAT heatid="23000" number="0" />
                <HEAT heatid="23001" number="1" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="10" agemax="-1" agemin="12" name="offene Wertung">
                  <RANKINGS>
                    <RANKING place="1" resultid="1514" />
                    <RANKING place="2" resultid="1515" />
                    <RANKING place="4" resultid="1516" />
                    <RANKING place="3" resultid="1517" />
                    <RANKING place="5" resultid="1518" />
                    <RANKING place="6" resultid="1520" />
                    <RANKING place="7" resultid="1521" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11" agemax="-1" agemin="12" name="Internationale offene Wertung">
                  <RANKINGS>
                    <RANKING place="1" resultid="1514" />
                    <RANKING place="2" resultid="1515" />
                    <RANKING place="4" resultid="1516" />
                    <RANKING place="3" resultid="1517" />
                    <RANKING place="6" resultid="1518" />
                    <RANKING place="5" resultid="1519" />
                    <RANKING place="7" resultid="1520" />
                    <RANKING place="8" resultid="1521" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="24" number="110" gender="M" round="FIN">
              <SWIMSTYLE stroke="SURFACE" relaycount="1" distance="200" />
              <HEATS>
                <HEAT heatid="24000" number="0" />
                <HEAT heatid="24001" number="1" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="10" agemax="-1" agemin="12" name="offene Wertung">
                  <RANKINGS>
                    <RANKING place="1" resultid="1527" />
                    <RANKING place="2" resultid="1528" />
                    <RANKING place="4" resultid="1529" />
                    <RANKING place="3" resultid="1530" />
                    <RANKING place="5" resultid="1531" />
                    <RANKING place="6" resultid="1532" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="25" number="311" gender="F" round="FIN">
              <SWIMSTYLE stroke="SURFACE" relaycount="1" distance="800" />
              <FEE value="650" currency="EUR" />
              <HEATS>
                <HEAT heatid="25001" number="1" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="4" agemax="13" agemin="12" name="Kategorie D" />
                <AGEGROUP agegroupid="3" agemax="15" agemin="14" name="Kategorie C">
                  <RANKINGS>
                    <RANKING place="1" resultid="466" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2" agemax="17" agemin="16" name="Kategorie B">
                  <RANKINGS>
                    <RANKING place="1" resultid="936" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1" agemax="21" agemin="18" name="Junior:innen">
                  <RANKINGS>
                    <RANKING place="4" resultid="77" />
                    <RANKING place="2" resultid="867" />
                    <RANKING place="3" resultid="1129" />
                    <RANKING place="1" resultid="1134" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="34" agemin="29" name="Master A" />
                <AGEGROUP agegroupid="6" agemax="44" agemin="35" name="Master B" />
                <AGEGROUP agegroupid="7" agemax="54" agemin="45" name="Master C" />
                <AGEGROUP agegroupid="8" agemax="64" agemin="55" name="Master D" />
                <AGEGROUP agegroupid="9" agemax="-1" agemin="65" name="Master E" />
                <AGEGROUP agegroupid="10" agemax="-1" agemin="12" name="offene Wertung">
                  <RANKINGS>
                    <RANKING place="6" resultid="77" />
                    <RANKING place="5" resultid="466" />
                    <RANKING place="3" resultid="867" />
                    <RANKING place="2" resultid="936" />
                    <RANKING place="4" resultid="1129" />
                    <RANKING place="1" resultid="1134" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11" agemax="-1" agemin="12" name="Internationale offene Wertung">
                  <RANKINGS>
                    <RANKING place="7" resultid="77" />
                    <RANKING place="3" resultid="172" />
                    <RANKING place="6" resultid="466" />
                    <RANKING place="4" resultid="867" />
                    <RANKING place="2" resultid="936" />
                    <RANKING place="5" resultid="1129" />
                    <RANKING place="1" resultid="1134" />
                    <RANKING place="8" resultid="1160" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="26" number="312" gender="M" round="FIN">
              <SWIMSTYLE stroke="SURFACE" relaycount="1" distance="800" />
              <FEE value="650" currency="EUR" />
              <HEATS>
                <HEAT heatid="26001" number="1" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="4" agemax="13" agemin="12" name="Kategorie D" />
                <AGEGROUP agegroupid="3" agemax="15" agemin="14" name="Kategorie C">
                  <RANKINGS>
                    <RANKING place="1" resultid="417" />
                    <RANKING place="2" resultid="450" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2" agemax="17" agemin="16" name="Kategorie B">
                  <RANKINGS>
                    <RANKING place="1" resultid="1177" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1" agemax="21" agemin="18" name="Junior:innen">
                  <RANKINGS>
                    <RANKING place="1" resultid="22" />
                    <RANKING place="2" resultid="388" />
                    <RANKING place="3" resultid="1347" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="34" agemin="29" name="Master A" />
                <AGEGROUP agegroupid="6" agemax="44" agemin="35" name="Master B" />
                <AGEGROUP agegroupid="7" agemax="54" agemin="45" name="Master C" />
                <AGEGROUP agegroupid="8" agemax="64" agemin="55" name="Master D" />
                <AGEGROUP agegroupid="9" agemax="-1" agemin="65" name="Master E" />
                <AGEGROUP agegroupid="10" agemax="-1" agemin="12" name="offene Wertung">
                  <RANKINGS>
                    <RANKING place="2" resultid="22" />
                    <RANKING place="3" resultid="388" />
                    <RANKING place="5" resultid="417" />
                    <RANKING place="7" resultid="450" />
                    <RANKING place="1" resultid="932" />
                    <RANKING place="6" resultid="1177" />
                    <RANKING place="4" resultid="1347" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11" agemax="-1" agemin="12" name="Internationale offene Wertung">
                  <RANKINGS>
                    <RANKING place="2" resultid="22" />
                    <RANKING place="5" resultid="218" />
                    <RANKING place="3" resultid="388" />
                    <RANKING place="6" resultid="417" />
                    <RANKING place="8" resultid="450" />
                    <RANKING place="1" resultid="932" />
                    <RANKING place="7" resultid="1177" />
                    <RANKING place="4" resultid="1347" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="27" number="313" gender="F" round="FIN">
              <SWIMSTYLE stroke="IMMERSION" technique="DIVE" relaycount="1" distance="400" />
              <FEE value="650" currency="EUR" />
              <HEATS>
                <HEAT heatid="27001" number="1" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="4" agemax="13" agemin="12" name="Kategorie D" />
                <AGEGROUP agegroupid="3" agemax="15" agemin="14" name="Kategorie C">
                  <RANKINGS>
                    <RANKING place="2" resultid="1030" />
                    <RANKING place="1" resultid="1232" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2" agemax="17" agemin="16" name="Kategorie B">
                  <RANKINGS>
                    <RANKING place="1" resultid="426" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1" agemax="21" agemin="18" name="Junior:innen">
                  <RANKINGS>
                    <RANKING place="1" resultid="768" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="34" agemin="29" name="Master A" />
                <AGEGROUP agegroupid="6" agemax="44" agemin="35" name="Master B" />
                <AGEGROUP agegroupid="7" agemax="54" agemin="45" name="Master C" />
                <AGEGROUP agegroupid="8" agemax="64" agemin="55" name="Master D" />
                <AGEGROUP agegroupid="9" agemax="-1" agemin="65" name="Master E" />
                <AGEGROUP agegroupid="10" agemax="-1" agemin="12" name="offene Wertung">
                  <RANKINGS>
                    <RANKING place="7" resultid="61" />
                    <RANKING place="5" resultid="72" />
                    <RANKING place="3" resultid="426" />
                    <RANKING place="6" resultid="768" />
                    <RANKING place="4" resultid="1030" />
                    <RANKING place="2" resultid="1232" />
                    <RANKING place="1" resultid="1302" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="28" number="314" gender="M" round="FIN">
              <SWIMSTYLE stroke="IMMERSION" technique="DIVE" relaycount="1" distance="400" />
              <FEE value="650" currency="EUR" />
              <HEATS>
                <HEAT heatid="28001" number="1" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="4" agemax="13" agemin="12" name="Kategorie D" />
                <AGEGROUP agegroupid="3" agemax="15" agemin="14" name="Kategorie C" />
                <AGEGROUP agegroupid="2" agemax="17" agemin="16" name="Kategorie B">
                  <RANKINGS>
                    <RANKING place="1" resultid="1178" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1" agemax="21" agemin="18" name="Junior:innen">
                  <RANKINGS>
                    <RANKING place="3" resultid="23" />
                    <RANKING place="5" resultid="160" />
                    <RANKING place="2" resultid="389" />
                    <RANKING place="1" resultid="476" />
                    <RANKING place="4" resultid="692" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="34" agemin="29" name="Master A" />
                <AGEGROUP agegroupid="6" agemax="44" agemin="35" name="Master B">
                  <RANKINGS>
                    <RANKING place="1" resultid="67" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7" agemax="54" agemin="45" name="Master C" />
                <AGEGROUP agegroupid="8" agemax="64" agemin="55" name="Master D" />
                <AGEGROUP agegroupid="9" agemax="-1" agemin="65" name="Master E" />
                <AGEGROUP agegroupid="10" agemax="-1" agemin="12" name="offene Wertung">
                  <RANKINGS>
                    <RANKING place="3" resultid="23" />
                    <RANKING place="6" resultid="67" />
                    <RANKING place="5" resultid="160" />
                    <RANKING place="2" resultid="389" />
                    <RANKING place="1" resultid="476" />
                    <RANKING place="4" resultid="692" />
                    <RANKING place="7" resultid="1178" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11" agemax="-1" agemin="12" name="Internationale offene Wertung">
                  <RANKINGS>
                    <RANKING place="4" resultid="23" />
                    <RANKING place="7" resultid="67" />
                    <RANKING place="6" resultid="160" />
                    <RANKING place="3" resultid="389" />
                    <RANKING place="2" resultid="476" />
                    <RANKING place="5" resultid="692" />
                    <RANKING place="1" resultid="1172" />
                    <RANKING place="8" resultid="1178" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="29" number="15" gender="X" round="TIM">
              <SWIMSTYLE stroke="SURFACE" relaycount="4" distance="50" />
              <FEE value="1000" currency="EUR" />
              <HEATS>
                <HEAT heatid="29001" number="1" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="5" agemax="-1" agemin="176" easy.ak="176" calculate="TOTAL" name="Master I" />
                <AGEGROUP agegroupid="6" agemax="-1" agemin="399" easy.ak="399" calculate="TOTAL" name="Master II">
                  <RANKINGS>
                    <RANKING place="2" resultid="1" />
                    <RANKING place="1" resultid="990" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="30" number="16" gender="X" round="TIM">
              <SWIMSTYLE stroke="SURFACE" relaycount="4" distance="50" />
              <FEE value="1000" currency="EUR" />
              <HEATS>
                <HEAT heatid="30001" number="1" />
                <HEAT heatid="30002" number="2" />
                <HEAT heatid="30003" number="3" />
                <HEAT heatid="30004" number="4" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="4" agemax="13" agemin="12" name="Kategorie D">
                  <RANKINGS>
                    <RANKING place="1" resultid="566" />
                    <RANKING place="2" resultid="1072" />
                    <RANKING place="3" resultid="1340" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3" agemax="15" agemin="14" name="Kategorie C">
                  <RANKINGS>
                    <RANKING place="1" resultid="410" />
                    <RANKING place="3" resultid="503" />
                    <RANKING place="4" resultid="568" />
                    <RANKING place="6" resultid="665" />
                    <RANKING place="5" resultid="819" />
                    <RANKING place="2" resultid="1185" />
                    <RANKING place="7" resultid="1341" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2" agemax="17" agemin="16" name="Kategorie B">
                  <RANKINGS>
                    <RANKING place="4" resultid="253" />
                    <RANKING place="2" resultid="910" />
                    <RANKING place="3" resultid="1079" />
                    <RANKING place="1" resultid="1116" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1" agemax="21" agemin="18" name="Junior:innen">
                  <RANKINGS>
                    <RANKING place="3" resultid="252" />
                    <RANKING place="1" resultid="408" />
                    <RANKING place="4" resultid="1186" />
                    <RANKING place="2" resultid="1328" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10" agemax="-1" agemin="12" name="offene Wertung">
                  <RANKINGS>
                    <RANKING place="15" resultid="91" />
                    <RANKING place="8" resultid="252" />
                    <RANKING place="12" resultid="253" />
                    <RANKING place="3" resultid="408" />
                    <RANKING place="10" resultid="410" />
                    <RANKING place="14" resultid="503" />
                    <RANKING place="19" resultid="566" />
                    <RANKING place="16" resultid="568" />
                    <RANKING place="18" resultid="665" />
                    <RANKING place="4" resultid="818" />
                    <RANKING place="17" resultid="819" />
                    <RANKING place="1" resultid="906" />
                    <RANKING place="7" resultid="910" />
                    <RANKING place="22" resultid="1072" />
                    <RANKING place="11" resultid="1079" />
                    <RANKING place="2" resultid="1113" />
                    <RANKING place="6" resultid="1116" />
                    <RANKING place="13" resultid="1185" />
                    <RANKING place="9" resultid="1186" />
                    <RANKING place="5" resultid="1328" />
                    <RANKING place="20" resultid="1338" />
                    <RANKING place="23" resultid="1340" />
                    <RANKING place="21" resultid="1341" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11" agemax="-1" agemin="12" name="Internationale offene Wertung">
                  <RANKINGS>
                    <RANKING place="16" resultid="91" />
                    <RANKING place="9" resultid="252" />
                    <RANKING place="13" resultid="253" />
                    <RANKING place="3" resultid="408" />
                    <RANKING place="11" resultid="410" />
                    <RANKING place="15" resultid="503" />
                    <RANKING place="20" resultid="566" />
                    <RANKING place="17" resultid="568" />
                    <RANKING place="19" resultid="665" />
                    <RANKING place="5" resultid="818" />
                    <RANKING place="18" resultid="819" />
                    <RANKING place="1" resultid="906" />
                    <RANKING place="8" resultid="910" />
                    <RANKING place="4" resultid="912" />
                    <RANKING place="23" resultid="1072" />
                    <RANKING place="12" resultid="1079" />
                    <RANKING place="2" resultid="1113" />
                    <RANKING place="7" resultid="1116" />
                    <RANKING place="14" resultid="1185" />
                    <RANKING place="10" resultid="1186" />
                    <RANKING place="6" resultid="1328" />
                    <RANKING place="21" resultid="1338" />
                    <RANKING place="24" resultid="1340" />
                    <RANKING place="22" resultid="1341" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
          </EVENTS>
        </SESSION>
        <SESSION number="4" date="2023-05-14" daytime="09:20" officialmeeting="08:45" warmupfrom="08:00">
          <EVENTS>
            <EVENT eventid="31" number="17" gender="F" round="PRE">
              <SWIMSTYLE stroke="SURFACE" relaycount="1" distance="100" />
              <FEE value="650" currency="EUR" />
              <HEATS>
                <HEAT heatid="31001" number="1" />
                <HEAT heatid="31002" number="2" />
                <HEAT heatid="31003" number="3" />
                <HEAT heatid="31004" number="4" />
                <HEAT heatid="31005" number="5" />
                <HEAT heatid="31006" number="6" />
                <HEAT heatid="31007" number="7" />
                <HEAT heatid="31008" number="8" />
                <HEAT heatid="31009" number="9" />
                <HEAT heatid="31010" number="10" />
                <HEAT heatid="31011" number="11" />
                <HEAT heatid="31012" number="12" />
                <HEAT heatid="31013" number="13" />
                <HEAT heatid="31014" number="14" />
                <HEAT heatid="31015" number="15" />
                <HEAT heatid="31016" number="16" />
                <HEAT heatid="31017" number="17" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="4" agemax="13" agemin="12" name="Kategorie D">
                  <RANKINGS>
                    <RANKING place="13" resultid="237" />
                    <RANKING place="5" resultid="242" />
                    <RANKING place="21" resultid="305" />
                    <RANKING place="3" resultid="363" />
                    <RANKING place="19" resultid="394" />
                    <RANKING place="10" resultid="422" />
                    <RANKING place="6" resultid="495" />
                    <RANKING place="1" resultid="573" />
                    <RANKING place="14" resultid="670" />
                    <RANKING place="9" resultid="699" />
                    <RANKING place="7" resultid="728" />
                    <RANKING place="18" resultid="789" />
                    <RANKING place="11" resultid="793" />
                    <RANKING place="2" resultid="825" />
                    <RANKING place="16" resultid="834" />
                    <RANKING place="4" resultid="874" />
                    <RANKING place="12" resultid="880" />
                    <RANKING place="17" resultid="945" />
                    <RANKING place="20" resultid="1057" />
                    <RANKING place="8" resultid="1076" />
                    <RANKING place="22" resultid="1239" />
                    <RANKING place="23" resultid="1243" />
                    <RANKING place="26" resultid="1258" />
                    <RANKING place="15" resultid="1274" />
                    <RANKING place="24" resultid="1289" />
                    <RANKING place="25" resultid="1312" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3" agemax="15" agemin="14" name="Kategorie C">
                  <RANKINGS>
                    <RANKING place="16" resultid="156" />
                    <RANKING place="25" resultid="226" />
                    <RANKING place="9" resultid="277" />
                    <RANKING place="7" resultid="282" />
                    <RANKING place="13" resultid="286" />
                    <RANKING place="19" resultid="314" />
                    <RANKING place="6" resultid="379" />
                    <RANKING place="21" resultid="413" />
                    <RANKING place="12" resultid="439" />
                    <RANKING place="24" resultid="447" />
                    <RANKING place="5" resultid="467" />
                    <RANKING place="15" resultid="490" />
                    <RANKING place="18" resultid="533" />
                    <RANKING place="8" resultid="588" />
                    <RANKING place="23" resultid="599" />
                    <RANKING place="11" resultid="642" />
                    <RANKING place="22" resultid="844" />
                    <RANKING place="4" resultid="954" />
                    <RANKING place="3" resultid="1031" />
                    <RANKING place="10" resultid="1207" />
                    <RANKING place="2" resultid="1212" />
                    <RANKING place="1" resultid="1233" />
                    <RANKING place="28" resultid="1251" />
                    <RANKING place="17" resultid="1270" />
                    <RANKING place="14" resultid="1285" />
                    <RANKING place="27" resultid="1316" />
                    <RANKING place="26" resultid="1358" />
                    <RANKING place="20" resultid="1366" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2" agemax="17" agemin="16" name="Kategorie B">
                  <RANKINGS>
                    <RANKING place="23" resultid="146" />
                    <RANKING place="3" resultid="427" />
                    <RANKING place="18" resultid="435" />
                    <RANKING place="5" resultid="444" />
                    <RANKING place="12" resultid="486" />
                    <RANKING place="20" resultid="519" />
                    <RANKING place="17" resultid="627" />
                    <RANKING place="11" resultid="900" />
                    <RANKING place="2" resultid="937" />
                    <RANKING place="21" resultid="958" />
                    <RANKING place="6" resultid="1050" />
                    <RANKING place="8" resultid="1098" />
                    <RANKING place="13" resultid="1103" />
                    <RANKING place="10" resultid="1141" />
                    <RANKING place="7" resultid="1149" />
                    <RANKING place="22" resultid="1153" />
                    <RANKING place="1" resultid="1167" />
                    <RANKING place="14" resultid="1193" />
                    <RANKING place="19" resultid="1226" />
                    <RANKING place="15" resultid="1255" />
                    <RANKING place="9" resultid="1310" />
                    <RANKING place="16" resultid="1319" />
                    <RANKING place="4" resultid="1344" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1" agemax="21" agemin="18" name="Junior:innen">
                  <RANKINGS>
                    <RANKING place="8" resultid="78" />
                    <RANKING place="18" resultid="110" />
                    <RANKING place="4" resultid="247" />
                    <RANKING place="13" resultid="259" />
                    <RANKING place="9" resultid="296" />
                    <RANKING place="15" resultid="455" />
                    <RANKING place="11" resultid="536" />
                    <RANKING place="6" resultid="761" />
                    <RANKING place="7" resultid="769" />
                    <RANKING place="5" resultid="868" />
                    <RANKING place="16" resultid="884" />
                    <RANKING place="1" resultid="976" />
                    <RANKING place="17" resultid="1035" />
                    <RANKING place="14" resultid="1064" />
                    <RANKING place="10" resultid="1130" />
                    <RANKING place="3" resultid="1135" />
                    <RANKING place="2" resultid="1145" />
                    <RANKING place="19" resultid="1181" />
                    <RANKING place="12" resultid="1381" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="34" agemin="29" name="Master A">
                  <RANKINGS>
                    <RANKING place="1" resultid="7" />
                    <RANKING place="2" resultid="49" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6" agemax="44" agemin="35" name="Master B">
                  <RANKINGS>
                    <RANKING place="2" resultid="650" />
                    <RANKING place="3" resultid="775" />
                    <RANKING place="4" resultid="894" />
                    <RANKING place="1" resultid="997" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7" agemax="54" agemin="45" name="Master C">
                  <RANKINGS>
                    <RANKING place="2" resultid="839" />
                    <RANKING place="1" resultid="1020" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8" agemax="64" agemin="55" name="Master D">
                  <RANKINGS>
                    <RANKING place="1" resultid="659" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9" agemax="-1" agemin="65" name="Master E">
                  <RANKINGS>
                    <RANKING place="1" resultid="993" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10" agemax="-1" agemin="12" name="offene Wertung">
                  <RANKINGS>
                    <RANKING place="44" resultid="7" />
                    <RANKING place="103" resultid="49" />
                    <RANKING place="35" resultid="62" />
                    <RANKING place="33" resultid="73" />
                    <RANKING place="16" resultid="78" />
                    <RANKING place="19" resultid="85" />
                    <RANKING place="54" resultid="110" />
                    <RANKING place="65" resultid="119" />
                    <RANKING place="52" resultid="143" />
                    <RANKING place="88" resultid="146" />
                    <RANKING place="76" resultid="156" />
                    <RANKING place="102" resultid="226" />
                    <RANKING place="95" resultid="237" />
                    <RANKING place="75" resultid="242" />
                    <RANKING place="6" resultid="247" />
                    <RANKING place="29" resultid="259" />
                    <RANKING place="49" resultid="277" />
                    <RANKING place="45" resultid="282" />
                    <RANKING place="64" resultid="286" />
                    <RANKING place="56" resultid="291" />
                    <RANKING place="20" resultid="296" />
                    <RANKING place="110" resultid="305" />
                    <RANKING place="82" resultid="314" />
                    <RANKING place="60" resultid="363" />
                    <RANKING place="37" resultid="379" />
                    <RANKING place="105" resultid="394" />
                    <RANKING place="85" resultid="413" />
                    <RANKING place="90" resultid="422" />
                    <RANKING place="10" resultid="427" />
                    <RANKING place="58" resultid="435" />
                    <RANKING place="61" resultid="439" />
                    <RANKING place="15" resultid="444" />
                    <RANKING place="94" resultid="447" />
                    <RANKING place="47" resultid="455" />
                    <RANKING place="32" resultid="467" />
                    <RANKING place="39" resultid="486" />
                    <RANKING place="74" resultid="490" />
                    <RANKING place="80" resultid="495" />
                    <RANKING place="66" resultid="519" />
                    <RANKING place="78" resultid="533" />
                    <RANKING place="23" resultid="536" />
                    <RANKING place="43" resultid="573" />
                    <RANKING place="46" resultid="588" />
                    <RANKING place="92" resultid="599" />
                    <RANKING place="55" resultid="627" />
                    <RANKING place="59" resultid="642" />
                    <RANKING place="72" resultid="650" />
                    <RANKING place="112" resultid="659" />
                    <RANKING place="97" resultid="670" />
                    <RANKING place="89" resultid="699" />
                    <RANKING place="81" resultid="728" />
                    <RANKING place="11" resultid="761" />
                    <RANKING place="14" resultid="769" />
                    <RANKING place="96" resultid="775" />
                    <RANKING place="3" resultid="780" />
                    <RANKING place="101" resultid="789" />
                    <RANKING place="91" resultid="793" />
                    <RANKING place="57" resultid="825" />
                    <RANKING place="99" resultid="834" />
                    <RANKING place="79" resultid="839" />
                    <RANKING place="87" resultid="844" />
                    <RANKING place="8" resultid="868" />
                    <RANKING place="69" resultid="874" />
                    <RANKING place="93" resultid="880" />
                    <RANKING place="51" resultid="884" />
                    <RANKING place="109" resultid="894" />
                    <RANKING place="38" resultid="900" />
                    <RANKING place="31" resultid="920" />
                    <RANKING place="18" resultid="929" />
                    <RANKING place="9" resultid="937" />
                    <RANKING place="100" resultid="945" />
                    <RANKING place="30" resultid="954" />
                    <RANKING place="71" resultid="958" />
                    <RANKING place="1" resultid="976" />
                    <RANKING place="12" resultid="988" />
                    <RANKING place="116" resultid="993" />
                    <RANKING place="70" resultid="997" />
                    <RANKING place="67" resultid="1020" />
                    <RANKING place="28" resultid="1031" />
                    <RANKING place="53" resultid="1035" />
                    <RANKING place="17" resultid="1050" />
                    <RANKING place="106" resultid="1057" />
                    <RANKING place="36" resultid="1064" />
                    <RANKING place="84" resultid="1076" />
                    <RANKING place="24" resultid="1098" />
                    <RANKING place="40" resultid="1103" />
                    <RANKING place="22" resultid="1130" />
                    <RANKING place="5" resultid="1135" />
                    <RANKING place="34" resultid="1141" />
                    <RANKING place="2" resultid="1145" />
                    <RANKING place="21" resultid="1149" />
                    <RANKING place="86" resultid="1153" />
                    <RANKING place="63" resultid="1157" />
                    <RANKING place="4" resultid="1167" />
                    <RANKING place="68" resultid="1181" />
                    <RANKING place="41" resultid="1193" />
                    <RANKING place="50" resultid="1207" />
                    <RANKING place="25" resultid="1212" />
                    <RANKING place="62" resultid="1226" />
                    <RANKING place="7" resultid="1233" />
                    <RANKING place="111" resultid="1239" />
                    <RANKING place="113" resultid="1243" />
                    <RANKING place="108" resultid="1251" />
                    <RANKING place="42" resultid="1255" />
                    <RANKING place="117" resultid="1258" />
                    <RANKING place="77" resultid="1270" />
                    <RANKING place="98" resultid="1274" />
                    <RANKING place="73" resultid="1285" />
                    <RANKING place="114" resultid="1289" />
                    <RANKING place="26" resultid="1310" />
                    <RANKING place="115" resultid="1312" />
                    <RANKING place="107" resultid="1316" />
                    <RANKING place="48" resultid="1319" />
                    <RANKING place="13" resultid="1344" />
                    <RANKING place="104" resultid="1358" />
                    <RANKING place="83" resultid="1366" />
                    <RANKING place="27" resultid="1381" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11" agemax="-1" agemin="12" name="Internationale Wertung">
                  <RANKINGS>
                    <RANKING place="47" resultid="7" />
                    <RANKING place="55" resultid="43" />
                    <RANKING place="111" resultid="49" />
                    <RANKING place="37" resultid="62" />
                    <RANKING place="35" resultid="73" />
                    <RANKING place="17" resultid="78" />
                    <RANKING place="21" resultid="85" />
                    <RANKING place="58" resultid="110" />
                    <RANKING place="70" resultid="119" />
                    <RANKING place="56" resultid="143" />
                    <RANKING place="96" resultid="146" />
                    <RANKING place="81" resultid="156" />
                    <RANKING place="89" resultid="215" />
                    <RANKING place="110" resultid="226" />
                    <RANKING place="103" resultid="237" />
                    <RANKING place="80" resultid="242" />
                    <RANKING place="6" resultid="247" />
                    <RANKING place="31" resultid="259" />
                    <RANKING place="52" resultid="277" />
                    <RANKING place="48" resultid="282" />
                    <RANKING place="69" resultid="286" />
                    <RANKING place="60" resultid="291" />
                    <RANKING place="22" resultid="296" />
                    <RANKING place="118" resultid="305" />
                    <RANKING place="87" resultid="314" />
                    <RANKING place="64" resultid="363" />
                    <RANKING place="39" resultid="379" />
                    <RANKING place="113" resultid="394" />
                    <RANKING place="93" resultid="413" />
                    <RANKING place="98" resultid="422" />
                    <RANKING place="11" resultid="427" />
                    <RANKING place="62" resultid="435" />
                    <RANKING place="65" resultid="439" />
                    <RANKING place="16" resultid="444" />
                    <RANKING place="102" resultid="447" />
                    <RANKING place="50" resultid="455" />
                    <RANKING place="90" resultid="461" />
                    <RANKING place="34" resultid="467" />
                    <RANKING place="42" resultid="486" />
                    <RANKING place="79" resultid="490" />
                    <RANKING place="85" resultid="495" />
                    <RANKING place="71" resultid="519" />
                    <RANKING place="83" resultid="533" />
                    <RANKING place="25" resultid="536" />
                    <RANKING place="46" resultid="573" />
                    <RANKING place="49" resultid="588" />
                    <RANKING place="100" resultid="599" />
                    <RANKING place="59" resultid="627" />
                    <RANKING place="63" resultid="642" />
                    <RANKING place="77" resultid="650" />
                    <RANKING place="120" resultid="659" />
                    <RANKING place="105" resultid="670" />
                    <RANKING place="97" resultid="699" />
                    <RANKING place="68" resultid="709" />
                    <RANKING place="86" resultid="728" />
                    <RANKING place="12" resultid="761" />
                    <RANKING place="15" resultid="769" />
                    <RANKING place="104" resultid="775" />
                    <RANKING place="3" resultid="780" />
                    <RANKING place="109" resultid="789" />
                    <RANKING place="99" resultid="793" />
                    <RANKING place="61" resultid="825" />
                    <RANKING place="107" resultid="834" />
                    <RANKING place="84" resultid="839" />
                    <RANKING place="95" resultid="844" />
                    <RANKING place="9" resultid="868" />
                    <RANKING place="74" resultid="874" />
                    <RANKING place="101" resultid="880" />
                    <RANKING place="54" resultid="884" />
                    <RANKING place="117" resultid="894" />
                    <RANKING place="41" resultid="900" />
                    <RANKING place="33" resultid="920" />
                    <RANKING place="20" resultid="929" />
                    <RANKING place="10" resultid="937" />
                    <RANKING place="108" resultid="945" />
                    <RANKING place="32" resultid="954" />
                    <RANKING place="76" resultid="958" />
                    <RANKING place="7" resultid="963" />
                    <RANKING place="1" resultid="976" />
                    <RANKING place="92" resultid="980" />
                    <RANKING place="40" resultid="985" />
                    <RANKING place="13" resultid="988" />
                    <RANKING place="124" resultid="993" />
                    <RANKING place="75" resultid="997" />
                    <RANKING place="72" resultid="1020" />
                    <RANKING place="30" resultid="1031" />
                    <RANKING place="57" resultid="1035" />
                    <RANKING place="19" resultid="1050" />
                    <RANKING place="114" resultid="1057" />
                    <RANKING place="38" resultid="1064" />
                    <RANKING place="91" resultid="1076" />
                    <RANKING place="26" resultid="1098" />
                    <RANKING place="43" resultid="1103" />
                    <RANKING place="24" resultid="1130" />
                    <RANKING place="5" resultid="1135" />
                    <RANKING place="36" resultid="1141" />
                    <RANKING place="2" resultid="1145" />
                    <RANKING place="23" resultid="1149" />
                    <RANKING place="94" resultid="1153" />
                    <RANKING place="67" resultid="1157" />
                    <RANKING place="18" resultid="1161" />
                    <RANKING place="4" resultid="1167" />
                    <RANKING place="73" resultid="1181" />
                    <RANKING place="44" resultid="1193" />
                    <RANKING place="53" resultid="1207" />
                    <RANKING place="27" resultid="1212" />
                    <RANKING place="66" resultid="1226" />
                    <RANKING place="8" resultid="1233" />
                    <RANKING place="119" resultid="1239" />
                    <RANKING place="121" resultid="1243" />
                    <RANKING place="116" resultid="1251" />
                    <RANKING place="45" resultid="1255" />
                    <RANKING place="125" resultid="1258" />
                    <RANKING place="82" resultid="1270" />
                    <RANKING place="106" resultid="1274" />
                    <RANKING place="78" resultid="1285" />
                    <RANKING place="122" resultid="1289" />
                    <RANKING place="28" resultid="1310" />
                    <RANKING place="123" resultid="1312" />
                    <RANKING place="115" resultid="1316" />
                    <RANKING place="51" resultid="1319" />
                    <RANKING place="14" resultid="1344" />
                    <RANKING place="112" resultid="1358" />
                    <RANKING place="88" resultid="1366" />
                    <RANKING place="29" resultid="1381" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="32" number="18" gender="M" round="PRE">
              <SWIMSTYLE stroke="SURFACE" relaycount="1" distance="100" />
              <FEE value="650" currency="EUR" />
              <HEATS>
                <HEAT heatid="32001" number="1" />
                <HEAT heatid="32002" number="2" />
                <HEAT heatid="32003" number="3" />
                <HEAT heatid="32004" number="4" />
                <HEAT heatid="32005" number="5" />
                <HEAT heatid="32006" number="6" />
                <HEAT heatid="32007" number="7" />
                <HEAT heatid="32008" number="8" />
                <HEAT heatid="32009" number="9" />
                <HEAT heatid="32010" number="10" />
                <HEAT heatid="32011" number="11" />
                <HEAT heatid="32012" number="12" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="4" agemax="13" agemin="12" name="Kategorie D">
                  <RANKINGS>
                    <RANKING place="6" resultid="96" />
                    <RANKING place="3" resultid="270" />
                    <RANKING place="14" resultid="514" />
                    <RANKING place="12" resultid="592" />
                    <RANKING place="1" resultid="617" />
                    <RANKING place="4" resultid="622" />
                    <RANKING place="9" resultid="632" />
                    <RANKING place="5" resultid="676" />
                    <RANKING place="2" resultid="704" />
                    <RANKING place="8" resultid="733" />
                    <RANKING place="10" resultid="1091" />
                    <RANKING place="11" resultid="1094" />
                    <RANKING place="13" resultid="1189" />
                    <RANKING place="16" resultid="1247" />
                    <RANKING place="15" resultid="1300" />
                    <RANKING place="7" resultid="1306" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3" agemax="15" agemin="14" name="Kategorie C">
                  <RANKINGS>
                    <RANKING place="14" resultid="114" />
                    <RANKING place="11" resultid="130" />
                    <RANKING place="9" resultid="400" />
                    <RANKING place="5" resultid="451" />
                    <RANKING place="2" resultid="529" />
                    <RANKING place="6" resultid="602" />
                    <RANKING place="13" resultid="607" />
                    <RANKING place="3" resultid="718" />
                    <RANKING place="12" resultid="850" />
                    <RANKING place="15" resultid="857" />
                    <RANKING place="4" resultid="917" />
                    <RANKING place="8" resultid="1087" />
                    <RANKING place="7" resultid="1198" />
                    <RANKING place="10" resultid="1218" />
                    <RANKING place="1" resultid="1353" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2" agemax="17" agemin="16" name="Kategorie B">
                  <RANKINGS>
                    <RANKING place="8" resultid="102" />
                    <RANKING place="7" resultid="264" />
                    <RANKING place="1" resultid="636" />
                    <RANKING place="10" resultid="686" />
                    <RANKING place="6" resultid="722" />
                    <RANKING place="2" resultid="798" />
                    <RANKING place="3" resultid="924" />
                    <RANKING place="5" resultid="1083" />
                    <RANKING place="4" resultid="1120" />
                    <RANKING place="9" resultid="1373" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1" agemax="21" agemin="18" name="Junior:innen">
                  <RANKINGS>
                    <RANKING place="4" resultid="24" />
                    <RANKING place="9" resultid="188" />
                    <RANKING place="14" resultid="301" />
                    <RANKING place="15" resultid="309" />
                    <RANKING place="7" resultid="318" />
                    <RANKING place="2" resultid="390" />
                    <RANKING place="8" resultid="431" />
                    <RANKING place="1" resultid="477" />
                    <RANKING place="11" resultid="679" />
                    <RANKING place="6" resultid="693" />
                    <RANKING place="13" resultid="712" />
                    <RANKING place="12" resultid="862" />
                    <RANKING place="5" resultid="1203" />
                    <RANKING place="10" resultid="1222" />
                    <RANKING place="3" resultid="1264" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="34" agemin="29" name="Master A">
                  <RANKINGS>
                    <RANKING place="1" resultid="968" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6" agemax="44" agemin="35" name="Master B">
                  <RANKINGS>
                    <RANKING place="2" resultid="35" />
                    <RANKING place="1" resultid="68" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7" agemax="54" agemin="45" name="Master C">
                  <RANKINGS>
                    <RANKING place="1" resultid="183" />
                    <RANKING place="5" resultid="541" />
                    <RANKING place="2" resultid="611" />
                    <RANKING place="7" resultid="645" />
                    <RANKING place="3" resultid="892" />
                    <RANKING place="4" resultid="1004" />
                    <RANKING place="6" resultid="1015" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8" agemax="64" agemin="55" name="Master D">
                  <RANKINGS>
                    <RANKING place="1" resultid="14" />
                    <RANKING place="2" resultid="203" />
                    <RANKING place="3" resultid="480" />
                    <RANKING place="4" resultid="739" />
                    <RANKING place="5" resultid="829" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9" agemax="-1" agemin="65" name="Master E">
                  <RANKINGS>
                    <RANKING place="1" resultid="195" />
                    <RANKING place="3" resultid="755" />
                    <RANKING place="2" resultid="1321" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10" agemax="-1" agemin="12" name="offene Wertung">
                  <RANKINGS>
                    <RANKING place="39" resultid="14" />
                    <RANKING place="13" resultid="24" />
                    <RANKING place="43" resultid="35" />
                    <RANKING place="29" resultid="68" />
                    <RANKING place="63" resultid="96" />
                    <RANKING place="34" resultid="102" />
                    <RANKING place="61" resultid="114" />
                    <RANKING place="55" resultid="130" />
                    <RANKING place="38" resultid="183" />
                    <RANKING place="22" resultid="188" />
                    <RANKING place="64" resultid="195" />
                    <RANKING place="45" resultid="203" />
                    <RANKING place="27" resultid="264" />
                    <RANKING place="57" resultid="270" />
                    <RANKING place="33" resultid="301" />
                    <RANKING place="44" resultid="309" />
                    <RANKING place="18" resultid="318" />
                    <RANKING place="6" resultid="390" />
                    <RANKING place="47" resultid="400" />
                    <RANKING place="19" resultid="431" />
                    <RANKING place="31" resultid="451" />
                    <RANKING place="5" resultid="477" />
                    <RANKING place="49" resultid="480" />
                    <RANKING place="76" resultid="514" />
                    <RANKING place="20" resultid="529" />
                    <RANKING place="51" resultid="541" />
                    <RANKING place="14" resultid="558" />
                    <RANKING place="73" resultid="592" />
                    <RANKING place="35" resultid="602" />
                    <RANKING place="59" resultid="607" />
                    <RANKING place="41" resultid="611" />
                    <RANKING place="48" resultid="617" />
                    <RANKING place="60" resultid="622" />
                    <RANKING place="69" resultid="632" />
                    <RANKING place="2" resultid="636" />
                    <RANKING place="58" resultid="645" />
                    <RANKING place="62" resultid="676" />
                    <RANKING place="24" resultid="679" />
                    <RANKING place="42" resultid="686" />
                    <RANKING place="17" resultid="693" />
                    <RANKING place="53" resultid="704" />
                    <RANKING place="32" resultid="712" />
                    <RANKING place="21" resultid="718" />
                    <RANKING place="26" resultid="722" />
                    <RANKING place="67" resultid="733" />
                    <RANKING place="66" resultid="739" />
                    <RANKING place="78" resultid="755" />
                    <RANKING place="7" resultid="798" />
                    <RANKING place="70" resultid="829" />
                    <RANKING place="56" resultid="850" />
                    <RANKING place="68" resultid="857" />
                    <RANKING place="30" resultid="862" />
                    <RANKING place="46" resultid="892" />
                    <RANKING place="28" resultid="917" />
                    <RANKING place="11" resultid="924" />
                    <RANKING place="12" resultid="941" />
                    <RANKING place="1" resultid="948" />
                    <RANKING place="3" resultid="968" />
                    <RANKING place="50" resultid="1004" />
                    <RANKING place="54" resultid="1015" />
                    <RANKING place="25" resultid="1083" />
                    <RANKING place="40" resultid="1087" />
                    <RANKING place="71" resultid="1091" />
                    <RANKING place="72" resultid="1094" />
                    <RANKING place="16" resultid="1120" />
                    <RANKING place="9" resultid="1124" />
                    <RANKING place="74" resultid="1189" />
                    <RANKING place="36" resultid="1198" />
                    <RANKING place="15" resultid="1203" />
                    <RANKING place="52" resultid="1218" />
                    <RANKING place="23" resultid="1222" />
                    <RANKING place="79" resultid="1247" />
                    <RANKING place="8" resultid="1264" />
                    <RANKING place="77" resultid="1300" />
                    <RANKING place="65" resultid="1306" />
                    <RANKING place="75" resultid="1321" />
                    <RANKING place="10" resultid="1353" />
                    <RANKING place="4" resultid="1361" />
                    <RANKING place="37" resultid="1373" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11" agemax="-1" agemin="12" name="Internationale offene Wertung">
                  <RANKINGS>
                    <RANKING place="45" resultid="14" />
                    <RANKING place="13" resultid="24" />
                    <RANKING place="49" resultid="35" />
                    <RANKING place="34" resultid="68" />
                    <RANKING place="69" resultid="96" />
                    <RANKING place="39" resultid="102" />
                    <RANKING place="67" resultid="114" />
                    <RANKING place="61" resultid="130" />
                    <RANKING place="15" resultid="164" />
                    <RANKING place="16" resultid="168" />
                    <RANKING place="43" resultid="183" />
                    <RANKING place="26" resultid="188" />
                    <RANKING place="70" resultid="195" />
                    <RANKING place="51" resultid="203" />
                    <RANKING place="44" resultid="209" />
                    <RANKING place="24" resultid="219" />
                    <RANKING place="31" resultid="264" />
                    <RANKING place="63" resultid="270" />
                    <RANKING place="38" resultid="301" />
                    <RANKING place="50" resultid="309" />
                    <RANKING place="21" resultid="318" />
                    <RANKING place="6" resultid="390" />
                    <RANKING place="53" resultid="400" />
                    <RANKING place="22" resultid="431" />
                    <RANKING place="36" resultid="451" />
                    <RANKING place="5" resultid="477" />
                    <RANKING place="55" resultid="480" />
                    <RANKING place="82" resultid="514" />
                    <RANKING place="23" resultid="529" />
                    <RANKING place="57" resultid="541" />
                    <RANKING place="17" resultid="558" />
                    <RANKING place="79" resultid="592" />
                    <RANKING place="40" resultid="602" />
                    <RANKING place="65" resultid="607" />
                    <RANKING place="47" resultid="611" />
                    <RANKING place="54" resultid="617" />
                    <RANKING place="66" resultid="622" />
                    <RANKING place="75" resultid="632" />
                    <RANKING place="2" resultid="636" />
                    <RANKING place="64" resultid="645" />
                    <RANKING place="68" resultid="676" />
                    <RANKING place="28" resultid="679" />
                    <RANKING place="48" resultid="686" />
                    <RANKING place="20" resultid="693" />
                    <RANKING place="59" resultid="704" />
                    <RANKING place="37" resultid="712" />
                    <RANKING place="25" resultid="718" />
                    <RANKING place="30" resultid="722" />
                    <RANKING place="73" resultid="733" />
                    <RANKING place="72" resultid="739" />
                    <RANKING place="84" resultid="755" />
                    <RANKING place="7" resultid="798" />
                    <RANKING place="76" resultid="829" />
                    <RANKING place="62" resultid="850" />
                    <RANKING place="74" resultid="857" />
                    <RANKING place="35" resultid="862" />
                    <RANKING place="52" resultid="892" />
                    <RANKING place="32" resultid="917" />
                    <RANKING place="11" resultid="924" />
                    <RANKING place="12" resultid="941" />
                    <RANKING place="1" resultid="948" />
                    <RANKING place="3" resultid="968" />
                    <RANKING place="33" resultid="971" />
                    <RANKING place="56" resultid="1004" />
                    <RANKING place="60" resultid="1015" />
                    <RANKING place="29" resultid="1083" />
                    <RANKING place="46" resultid="1087" />
                    <RANKING place="77" resultid="1091" />
                    <RANKING place="78" resultid="1094" />
                    <RANKING place="19" resultid="1120" />
                    <RANKING place="9" resultid="1124" />
                    <RANKING place="14" resultid="1173" />
                    <RANKING place="80" resultid="1189" />
                    <RANKING place="41" resultid="1198" />
                    <RANKING place="18" resultid="1203" />
                    <RANKING place="58" resultid="1218" />
                    <RANKING place="27" resultid="1222" />
                    <RANKING place="85" resultid="1247" />
                    <RANKING place="8" resultid="1264" />
                    <RANKING place="83" resultid="1300" />
                    <RANKING place="71" resultid="1306" />
                    <RANKING place="81" resultid="1321" />
                    <RANKING place="10" resultid="1353" />
                    <RANKING place="4" resultid="1361" />
                    <RANKING place="42" resultid="1373" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="33" number="19" gender="F" round="TIM">
              <SWIMSTYLE stroke="SURFACE" relaycount="1" distance="400" />
              <FEE value="650" currency="EUR" />
              <HEATS>
                <HEAT heatid="33001" number="1" />
                <HEAT heatid="33002" number="2" />
                <HEAT heatid="33003" number="3" />
                <HEAT heatid="33004" number="4" />
                <HEAT heatid="33005" number="5" />
                <HEAT heatid="33006" number="6" />
                <HEAT heatid="33007" number="7" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="4" agemax="13" agemin="12" name="Kategorie D">
                  <RANKINGS>
                    <RANKING place="2" resultid="423" />
                    <RANKING place="10" resultid="548" />
                    <RANKING place="6" resultid="671" />
                    <RANKING place="9" resultid="790" />
                    <RANKING place="5" resultid="794" />
                    <RANKING place="1" resultid="826" />
                    <RANKING place="4" resultid="881" />
                    <RANKING place="8" resultid="1058" />
                    <RANKING place="3" resultid="1275" />
                    <RANKING place="7" resultid="1297" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3" agemax="15" agemin="14" name="Kategorie C">
                  <RANKINGS>
                    <RANKING place="12" resultid="227" />
                    <RANKING place="3" resultid="278" />
                    <RANKING place="8" resultid="414" />
                    <RANKING place="2" resultid="440" />
                    <RANKING place="1" resultid="468" />
                    <RANKING place="7" resultid="643" />
                    <RANKING place="10" resultid="845" />
                    <RANKING place="6" resultid="1208" />
                    <RANKING place="9" resultid="1278" />
                    <RANKING place="4" resultid="1286" />
                    <RANKING place="11" resultid="1317" />
                    <RANKING place="5" resultid="1367" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2" agemax="17" agemin="16" name="Kategorie B">
                  <RANKINGS>
                    <RANKING place="2" resultid="231" />
                    <RANKING place="4" resultid="384" />
                    <RANKING place="6" resultid="628" />
                    <RANKING place="7" resultid="901" />
                    <RANKING place="1" resultid="1104" />
                    <RANKING place="8" resultid="1154" />
                    <RANKING place="5" resultid="1194" />
                    <RANKING place="3" resultid="1256" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1" agemax="21" agemin="18" name="Junior:innen">
                  <RANKINGS>
                    <RANKING place="1" resultid="79" />
                    <RANKING place="5" resultid="111" />
                    <RANKING place="4" resultid="151" />
                    <RANKING place="2" resultid="537" />
                    <RANKING place="3" resultid="1131" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="34" agemin="29" name="Master A">
                  <RANKINGS>
                    <RANKING place="1" resultid="8" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6" agemax="44" agemin="35" name="Master B">
                  <RANKINGS>
                    <RANKING place="1" resultid="651" />
                    <RANKING place="2" resultid="776" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7" agemax="54" agemin="45" name="Master C">
                  <RANKINGS>
                    <RANKING place="1" resultid="30" />
                    <RANKING place="2" resultid="840" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8" agemax="64" agemin="55" name="Master D">
                  <RANKINGS>
                    <RANKING place="1" resultid="660" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9" agemax="-1" agemin="65" name="Master E" />
                <AGEGROUP agegroupid="10" agemax="-1" agemin="12" name="offene Wertung">
                  <RANKINGS>
                    <RANKING place="10" resultid="8" />
                    <RANKING place="14" resultid="30" />
                    <RANKING place="3" resultid="63" />
                    <RANKING place="4" resultid="79" />
                    <RANKING place="1" resultid="86" />
                    <RANKING place="12" resultid="111" />
                    <RANKING place="18" resultid="120" />
                    <RANKING place="9" resultid="151" />
                    <RANKING place="40" resultid="227" />
                    <RANKING place="8" resultid="231" />
                    <RANKING place="19" resultid="278" />
                    <RANKING place="13" resultid="384" />
                    <RANKING place="29" resultid="414" />
                    <RANKING place="23" resultid="423" />
                    <RANKING place="15" resultid="440" />
                    <RANKING place="2" resultid="468" />
                    <RANKING place="5" resultid="537" />
                    <RANKING place="43" resultid="548" />
                    <RANKING place="17" resultid="628" />
                    <RANKING place="28" resultid="643" />
                    <RANKING place="24" resultid="651" />
                    <RANKING place="44" resultid="660" />
                    <RANKING place="37" resultid="671" />
                    <RANKING place="34" resultid="776" />
                    <RANKING place="42" resultid="790" />
                    <RANKING place="35" resultid="794" />
                    <RANKING place="22" resultid="826" />
                    <RANKING place="27" resultid="840" />
                    <RANKING place="32" resultid="845" />
                    <RANKING place="33" resultid="881" />
                    <RANKING place="20" resultid="901" />
                    <RANKING place="41" resultid="1058" />
                    <RANKING place="7" resultid="1104" />
                    <RANKING place="6" resultid="1131" />
                    <RANKING place="36" resultid="1154" />
                    <RANKING place="16" resultid="1194" />
                    <RANKING place="26" resultid="1208" />
                    <RANKING place="11" resultid="1256" />
                    <RANKING place="31" resultid="1275" />
                    <RANKING place="30" resultid="1278" />
                    <RANKING place="21" resultid="1286" />
                    <RANKING place="39" resultid="1297" />
                    <RANKING place="38" resultid="1317" />
                    <RANKING place="25" resultid="1367" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11" agemax="-1" agemin="12" name="Internationale offene Wertung">
                  <RANKINGS>
                    <RANKING place="11" resultid="8" />
                    <RANKING place="17" resultid="30" />
                    <RANKING place="15" resultid="44" />
                    <RANKING place="3" resultid="63" />
                    <RANKING place="4" resultid="79" />
                    <RANKING place="1" resultid="86" />
                    <RANKING place="14" resultid="111" />
                    <RANKING place="21" resultid="120" />
                    <RANKING place="10" resultid="151" />
                    <RANKING place="44" resultid="227" />
                    <RANKING place="9" resultid="231" />
                    <RANKING place="23" resultid="278" />
                    <RANKING place="16" resultid="384" />
                    <RANKING place="33" resultid="414" />
                    <RANKING place="27" resultid="423" />
                    <RANKING place="18" resultid="440" />
                    <RANKING place="2" resultid="468" />
                    <RANKING place="5" resultid="537" />
                    <RANKING place="47" resultid="548" />
                    <RANKING place="12" resultid="579" />
                    <RANKING place="20" resultid="628" />
                    <RANKING place="32" resultid="643" />
                    <RANKING place="28" resultid="651" />
                    <RANKING place="48" resultid="660" />
                    <RANKING place="41" resultid="671" />
                    <RANKING place="22" resultid="710" />
                    <RANKING place="38" resultid="776" />
                    <RANKING place="46" resultid="790" />
                    <RANKING place="39" resultid="794" />
                    <RANKING place="26" resultid="826" />
                    <RANKING place="31" resultid="840" />
                    <RANKING place="36" resultid="845" />
                    <RANKING place="37" resultid="881" />
                    <RANKING place="24" resultid="901" />
                    <RANKING place="7" resultid="986" />
                    <RANKING place="45" resultid="1058" />
                    <RANKING place="8" resultid="1104" />
                    <RANKING place="6" resultid="1131" />
                    <RANKING place="40" resultid="1154" />
                    <RANKING place="19" resultid="1194" />
                    <RANKING place="30" resultid="1208" />
                    <RANKING place="13" resultid="1256" />
                    <RANKING place="35" resultid="1275" />
                    <RANKING place="34" resultid="1278" />
                    <RANKING place="25" resultid="1286" />
                    <RANKING place="43" resultid="1297" />
                    <RANKING place="42" resultid="1317" />
                    <RANKING place="29" resultid="1367" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="34" number="20" gender="M" round="TIM">
              <SWIMSTYLE stroke="SURFACE" relaycount="1" distance="400" />
              <FEE value="650" currency="EUR" />
              <HEATS>
                <HEAT heatid="34001" number="1" />
                <HEAT heatid="34002" number="2" />
                <HEAT heatid="34003" number="3" />
                <HEAT heatid="34004" number="4" />
                <HEAT heatid="34005" number="5" />
                <HEAT heatid="34006" number="6" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="4" agemax="13" agemin="12" name="Kategorie D">
                  <RANKINGS>
                    <RANKING place="4" resultid="97" />
                    <RANKING place="1" resultid="271" />
                    <RANKING place="9" resultid="515" />
                    <RANKING place="2" resultid="618" />
                    <RANKING place="5" resultid="623" />
                    <RANKING place="8" resultid="677" />
                    <RANKING place="3" resultid="705" />
                    <RANKING place="7" resultid="1190" />
                    <RANKING place="6" resultid="1307" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3" agemax="15" agemin="14" name="Kategorie C">
                  <RANKINGS>
                    <RANKING place="12" resultid="115" />
                    <RANKING place="10" resultid="131" />
                    <RANKING place="7" resultid="138" />
                    <RANKING place="8" resultid="401" />
                    <RANKING place="2" resultid="452" />
                    <RANKING place="11" resultid="510" />
                    <RANKING place="6" resultid="525" />
                    <RANKING place="13" resultid="696" />
                    <RANKING place="14" resultid="851" />
                    <RANKING place="1" resultid="918" />
                    <RANKING place="4" resultid="1088" />
                    <RANKING place="3" resultid="1199" />
                    <RANKING place="9" resultid="1219" />
                    <RANKING place="15" resultid="1292" />
                    <RANKING place="5" resultid="1325" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2" agemax="17" agemin="16" name="Kategorie B">
                  <RANKINGS>
                    <RANKING place="2" resultid="103" />
                    <RANKING place="1" resultid="1179" />
                    <RANKING place="3" resultid="1374" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1" agemax="21" agemin="18" name="Junior:innen">
                  <RANKINGS>
                    <RANKING place="2" resultid="161" />
                    <RANKING place="3" resultid="302" />
                    <RANKING place="4" resultid="310" />
                    <RANKING place="1" resultid="694" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="34" agemin="29" name="Master A" />
                <AGEGROUP agegroupid="6" agemax="44" agemin="35" name="Master B">
                  <RANKINGS>
                    <RANKING place="2" resultid="36" />
                    <RANKING place="1" resultid="69" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7" agemax="54" agemin="45" name="Master C">
                  <RANKINGS>
                    <RANKING place="2" resultid="802" />
                    <RANKING place="1" resultid="1011" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8" agemax="64" agemin="55" name="Master D">
                  <RANKINGS>
                    <RANKING place="1" resultid="15" />
                    <RANKING place="3" resultid="57" />
                    <RANKING place="4" resultid="740" />
                    <RANKING place="2" resultid="1025" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9" agemax="-1" agemin="65" name="Master E">
                  <RANKINGS>
                    <RANKING place="1" resultid="756" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10" agemax="-1" agemin="12" name="offene Wertung">
                  <RANKINGS>
                    <RANKING place="6" resultid="15" />
                    <RANKING place="18" resultid="36" />
                    <RANKING place="26" resultid="57" />
                    <RANKING place="10" resultid="69" />
                    <RANKING place="27" resultid="97" />
                    <RANKING place="11" resultid="103" />
                    <RANKING place="30" resultid="115" />
                    <RANKING place="25" resultid="131" />
                    <RANKING place="19" resultid="138" />
                    <RANKING place="2" resultid="161" />
                    <RANKING place="17" resultid="271" />
                    <RANKING place="12" resultid="302" />
                    <RANKING place="14" resultid="310" />
                    <RANKING place="21" resultid="401" />
                    <RANKING place="7" resultid="452" />
                    <RANKING place="28" resultid="510" />
                    <RANKING place="38" resultid="515" />
                    <RANKING place="16" resultid="525" />
                    <RANKING place="23" resultid="618" />
                    <RANKING place="29" resultid="623" />
                    <RANKING place="35" resultid="677" />
                    <RANKING place="1" resultid="694" />
                    <RANKING place="32" resultid="696" />
                    <RANKING place="24" resultid="705" />
                    <RANKING place="39" resultid="740" />
                    <RANKING place="40" resultid="756" />
                    <RANKING place="33" resultid="802" />
                    <RANKING place="36" resultid="851" />
                    <RANKING place="5" resultid="918" />
                    <RANKING place="4" resultid="1011" />
                    <RANKING place="20" resultid="1025" />
                    <RANKING place="9" resultid="1088" />
                    <RANKING place="3" resultid="1179" />
                    <RANKING place="34" resultid="1190" />
                    <RANKING place="8" resultid="1199" />
                    <RANKING place="22" resultid="1219" />
                    <RANKING place="37" resultid="1292" />
                    <RANKING place="31" resultid="1307" />
                    <RANKING place="15" resultid="1325" />
                    <RANKING place="13" resultid="1374" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11" agemax="-1" agemin="12" name="Internationale offene Wertung">
                  <RANKINGS>
                    <RANKING place="6" resultid="15" />
                    <RANKING place="18" resultid="36" />
                    <RANKING place="26" resultid="57" />
                    <RANKING place="10" resultid="69" />
                    <RANKING place="27" resultid="97" />
                    <RANKING place="11" resultid="103" />
                    <RANKING place="30" resultid="115" />
                    <RANKING place="25" resultid="131" />
                    <RANKING place="19" resultid="138" />
                    <RANKING place="2" resultid="161" />
                    <RANKING place="17" resultid="271" />
                    <RANKING place="12" resultid="302" />
                    <RANKING place="14" resultid="310" />
                    <RANKING place="21" resultid="401" />
                    <RANKING place="7" resultid="452" />
                    <RANKING place="28" resultid="510" />
                    <RANKING place="38" resultid="515" />
                    <RANKING place="16" resultid="525" />
                    <RANKING place="23" resultid="618" />
                    <RANKING place="29" resultid="623" />
                    <RANKING place="35" resultid="677" />
                    <RANKING place="1" resultid="694" />
                    <RANKING place="32" resultid="696" />
                    <RANKING place="24" resultid="705" />
                    <RANKING place="39" resultid="740" />
                    <RANKING place="40" resultid="756" />
                    <RANKING place="33" resultid="802" />
                    <RANKING place="36" resultid="851" />
                    <RANKING place="5" resultid="918" />
                    <RANKING place="4" resultid="1011" />
                    <RANKING place="20" resultid="1025" />
                    <RANKING place="9" resultid="1088" />
                    <RANKING place="3" resultid="1179" />
                    <RANKING place="34" resultid="1190" />
                    <RANKING place="8" resultid="1199" />
                    <RANKING place="22" resultid="1219" />
                    <RANKING place="37" resultid="1292" />
                    <RANKING place="31" resultid="1307" />
                    <RANKING place="15" resultid="1325" />
                    <RANKING place="13" resultid="1374" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="35" number="21" gender="F" round="TIM">
              <SWIMSTYLE stroke="IMMERSION" technique="DIVE" relaycount="1" distance="50" />
              <FEE value="650" currency="EUR" />
              <HEATS>
                <HEAT heatid="35001" number="1" />
                <HEAT heatid="35002" number="2" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="4" agemax="13" agemin="12" name="Kategorie D">
                  <RANKINGS>
                    <RANKING place="8" resultid="238" />
                    <RANKING place="6" resultid="243" />
                    <RANKING place="11" resultid="306" />
                    <RANKING place="3" resultid="364" />
                    <RANKING place="9" resultid="375" />
                    <RANKING place="2" resultid="496" />
                    <RANKING place="1" resultid="574" />
                    <RANKING place="7" resultid="700" />
                    <RANKING place="4" resultid="729" />
                    <RANKING place="9" resultid="1059" />
                    <RANKING place="5" resultid="1078" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="13" agemin="12" name="Internationale offene Wertung">
                  <RANKINGS>
                    <RANKING place="1" resultid="45" />
                    <RANKING place="10" resultid="238" />
                    <RANKING place="7" resultid="243" />
                    <RANKING place="13" resultid="306" />
                    <RANKING place="4" resultid="364" />
                    <RANKING place="11" resultid="375" />
                    <RANKING place="3" resultid="496" />
                    <RANKING place="2" resultid="574" />
                    <RANKING place="8" resultid="700" />
                    <RANKING place="5" resultid="729" />
                    <RANKING place="9" resultid="981" />
                    <RANKING place="11" resultid="1059" />
                    <RANKING place="6" resultid="1078" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="36" number="22" gender="M" round="TIM">
              <SWIMSTYLE stroke="IMMERSION" technique="DIVE" relaycount="1" distance="50" />
              <FEE value="650" currency="EUR" />
              <HEATS>
                <HEAT heatid="36001" number="1" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="4" agemax="13" agemin="12" name="Kategorie D">
                  <RANKINGS>
                    <RANKING place="2" resultid="272" />
                    <RANKING place="1" resultid="619" />
                    <RANKING place="4" resultid="678" />
                    <RANKING place="3" resultid="706" />
                    <RANKING place="5" resultid="734" />
                    <RANKING place="6" resultid="1248" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="37" number="23" gender="F" round="PRE">
              <SWIMSTYLE stroke="APNEA" relaycount="1" distance="50" />
              <FEE value="650" currency="EUR" />
              <HEATS>
                <HEAT heatid="37001" number="1" />
                <HEAT heatid="37002" number="2" />
                <HEAT heatid="37003" number="3" />
                <HEAT heatid="37004" number="4" />
                <HEAT heatid="37005" number="5" />
                <HEAT heatid="37006" number="6" />
                <HEAT heatid="37007" number="7" />
                <HEAT heatid="37008" number="8" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="3" agemax="15" agemin="14" name="Kategorie C">
                  <RANKINGS>
                    <RANKING place="10" resultid="279" />
                    <RANKING place="7" resultid="283" />
                    <RANKING place="13" resultid="315" />
                    <RANKING place="4" resultid="380" />
                    <RANKING place="5" resultid="469" />
                    <RANKING place="12" resultid="491" />
                    <RANKING place="9" resultid="589" />
                    <RANKING place="14" resultid="846" />
                    <RANKING place="3" resultid="955" />
                    <RANKING place="2" resultid="1032" />
                    <RANKING place="11" resultid="1209" />
                    <RANKING place="6" resultid="1213" />
                    <RANKING place="1" resultid="1234" />
                    <RANKING place="15" resultid="1252" />
                    <RANKING place="8" resultid="1271" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2" agemax="17" agemin="16" name="Kategorie B">
                  <RANKINGS>
                    <RANKING place="7" resultid="232" />
                    <RANKING place="17" resultid="385" />
                    <RANKING place="4" resultid="429" />
                    <RANKING place="12" resultid="436" />
                    <RANKING place="1" resultid="445" />
                    <RANKING place="11" resultid="487" />
                    <RANKING place="9" resultid="520" />
                    <RANKING place="15" resultid="629" />
                    <RANKING place="10" resultid="902" />
                    <RANKING place="16" resultid="959" />
                    <RANKING place="3" resultid="1051" />
                    <RANKING place="6" resultid="1099" />
                    <RANKING place="8" resultid="1142" />
                    <RANKING place="5" resultid="1150" />
                    <RANKING place="18" resultid="1155" />
                    <RANKING place="13" resultid="1195" />
                    <RANKING place="14" resultid="1228" />
                    <RANKING place="2" resultid="1345" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1" agemax="21" agemin="18" name="Junior:innen">
                  <RANKINGS>
                    <RANKING place="11" resultid="152" />
                    <RANKING place="1" resultid="248" />
                    <RANKING place="11" resultid="260" />
                    <RANKING place="7" resultid="297" />
                    <RANKING place="15" resultid="456" />
                    <RANKING place="9" resultid="538" />
                    <RANKING place="3" resultid="762" />
                    <RANKING place="6" resultid="771" />
                    <RANKING place="10" resultid="854" />
                    <RANKING place="5" resultid="870" />
                    <RANKING place="14" resultid="885" />
                    <RANKING place="13" resultid="1036" />
                    <RANKING place="8" resultid="1048" />
                    <RANKING place="2" resultid="1146" />
                    <RANKING place="16" resultid="1182" />
                    <RANKING place="4" resultid="1386" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="34" agemin="29" name="Master A" />
                <AGEGROUP agegroupid="6" agemax="44" agemin="35" name="Master B">
                  <RANKINGS>
                    <RANKING place="1" resultid="652" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7" agemax="54" agemin="45" name="Master C">
                  <RANKINGS>
                    <RANKING place="1" resultid="31" />
                    <RANKING place="2" resultid="1021" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8" agemax="64" agemin="55" name="Master D">
                  <RANKINGS>
                    <RANKING place="1" resultid="661" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9" agemax="-1" agemin="65" name="Master E" />
                <AGEGROUP agegroupid="10" agemax="-1" agemin="14" name="offene Wertung">
                  <RANKINGS>
                    <RANKING place="39" resultid="31" />
                    <RANKING place="23" resultid="74" />
                    <RANKING place="26" resultid="152" />
                    <RANKING place="24" resultid="232" />
                    <RANKING place="2" resultid="248" />
                    <RANKING place="26" resultid="260" />
                    <RANKING place="46" resultid="279" />
                    <RANKING place="34" resultid="283" />
                    <RANKING place="38" resultid="292" />
                    <RANKING place="15" resultid="297" />
                    <RANKING place="54" resultid="315" />
                    <RANKING place="22" resultid="380" />
                    <RANKING place="51" resultid="385" />
                    <RANKING place="12" resultid="429" />
                    <RANKING place="36" resultid="436" />
                    <RANKING place="3" resultid="445" />
                    <RANKING place="42" resultid="456" />
                    <RANKING place="28" resultid="469" />
                    <RANKING place="35" resultid="487" />
                    <RANKING place="52" resultid="491" />
                    <RANKING place="30" resultid="520" />
                    <RANKING place="20" resultid="538" />
                    <RANKING place="45" resultid="589" />
                    <RANKING place="44" resultid="629" />
                    <RANKING place="55" resultid="652" />
                    <RANKING place="58" resultid="661" />
                    <RANKING place="6" resultid="762" />
                    <RANKING place="14" resultid="771" />
                    <RANKING place="1" resultid="781" />
                    <RANKING place="56" resultid="846" />
                    <RANKING place="25" resultid="854" />
                    <RANKING place="10" resultid="870" />
                    <RANKING place="41" resultid="885" />
                    <RANKING place="31" resultid="902" />
                    <RANKING place="21" resultid="921" />
                    <RANKING place="18" resultid="955" />
                    <RANKING place="49" resultid="959" />
                    <RANKING place="9" resultid="989" />
                    <RANKING place="47" resultid="1021" />
                    <RANKING place="13" resultid="1032" />
                    <RANKING place="33" resultid="1036" />
                    <RANKING place="19" resultid="1048" />
                    <RANKING place="11" resultid="1051" />
                    <RANKING place="17" resultid="1099" />
                    <RANKING place="28" resultid="1142" />
                    <RANKING place="4" resultid="1146" />
                    <RANKING place="16" resultid="1150" />
                    <RANKING place="53" resultid="1155" />
                    <RANKING place="50" resultid="1182" />
                    <RANKING place="37" resultid="1195" />
                    <RANKING place="48" resultid="1209" />
                    <RANKING place="32" resultid="1213" />
                    <RANKING place="40" resultid="1228" />
                    <RANKING place="7" resultid="1234" />
                    <RANKING place="57" resultid="1252" />
                    <RANKING place="43" resultid="1271" />
                    <RANKING place="5" resultid="1345" />
                    <RANKING place="8" resultid="1386" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11" agemax="-1" agemin="14" name="Internationale offene Wertung">
                  <RANKINGS>
                    <RANKING place="41" resultid="31" />
                    <RANKING place="24" resultid="74" />
                    <RANKING place="27" resultid="152" />
                    <RANKING place="25" resultid="232" />
                    <RANKING place="3" resultid="248" />
                    <RANKING place="27" resultid="260" />
                    <RANKING place="48" resultid="279" />
                    <RANKING place="36" resultid="283" />
                    <RANKING place="40" resultid="292" />
                    <RANKING place="16" resultid="297" />
                    <RANKING place="56" resultid="315" />
                    <RANKING place="23" resultid="380" />
                    <RANKING place="53" resultid="385" />
                    <RANKING place="13" resultid="429" />
                    <RANKING place="38" resultid="436" />
                    <RANKING place="4" resultid="445" />
                    <RANKING place="44" resultid="456" />
                    <RANKING place="29" resultid="469" />
                    <RANKING place="37" resultid="487" />
                    <RANKING place="54" resultid="491" />
                    <RANKING place="31" resultid="520" />
                    <RANKING place="21" resultid="538" />
                    <RANKING place="35" resultid="580" />
                    <RANKING place="47" resultid="589" />
                    <RANKING place="46" resultid="629" />
                    <RANKING place="57" resultid="652" />
                    <RANKING place="60" resultid="661" />
                    <RANKING place="7" resultid="762" />
                    <RANKING place="15" resultid="771" />
                    <RANKING place="1" resultid="781" />
                    <RANKING place="58" resultid="846" />
                    <RANKING place="26" resultid="854" />
                    <RANKING place="11" resultid="870" />
                    <RANKING place="43" resultid="885" />
                    <RANKING place="32" resultid="902" />
                    <RANKING place="22" resultid="921" />
                    <RANKING place="19" resultid="955" />
                    <RANKING place="51" resultid="959" />
                    <RANKING place="2" resultid="964" />
                    <RANKING place="10" resultid="989" />
                    <RANKING place="49" resultid="1021" />
                    <RANKING place="14" resultid="1032" />
                    <RANKING place="34" resultid="1036" />
                    <RANKING place="20" resultid="1048" />
                    <RANKING place="12" resultid="1051" />
                    <RANKING place="18" resultid="1099" />
                    <RANKING place="29" resultid="1142" />
                    <RANKING place="5" resultid="1146" />
                    <RANKING place="17" resultid="1150" />
                    <RANKING place="55" resultid="1155" />
                    <RANKING place="52" resultid="1182" />
                    <RANKING place="39" resultid="1195" />
                    <RANKING place="50" resultid="1209" />
                    <RANKING place="33" resultid="1213" />
                    <RANKING place="42" resultid="1228" />
                    <RANKING place="8" resultid="1234" />
                    <RANKING place="59" resultid="1252" />
                    <RANKING place="45" resultid="1271" />
                    <RANKING place="6" resultid="1345" />
                    <RANKING place="9" resultid="1386" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="38" number="24" gender="M" round="PRE">
              <SWIMSTYLE stroke="APNEA" relaycount="1" distance="50" />
              <FEE value="650" currency="EUR" />
              <HEATS>
                <HEAT heatid="38001" number="1" />
                <HEAT heatid="38002" number="2" />
                <HEAT heatid="38003" number="3" />
                <HEAT heatid="38004" number="4" />
                <HEAT heatid="38005" number="5" />
                <HEAT heatid="38006" number="6" />
                <HEAT heatid="38007" number="7" />
                <HEAT heatid="38008" number="8" />
                <HEAT heatid="38009" number="9" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="3" agemax="15" agemin="14" name="Kategorie C">
                  <RANKINGS>
                    <RANKING place="13" resultid="132" />
                    <RANKING place="7" resultid="139" />
                    <RANKING place="14" resultid="402" />
                    <RANKING place="6" resultid="453" />
                    <RANKING place="11" resultid="511" />
                    <RANKING place="8" resultid="526" />
                    <RANKING place="2" resultid="530" />
                    <RANKING place="9" resultid="603" />
                    <RANKING place="15" resultid="682" />
                    <RANKING place="16" resultid="697" />
                    <RANKING place="1" resultid="719" />
                    <RANKING place="12" resultid="852" />
                    <RANKING place="4" resultid="919" />
                    <RANKING place="10" resultid="1107" />
                    <RANKING place="5" resultid="1200" />
                    <RANKING place="17" resultid="1293" />
                    <RANKING place="3" resultid="1354" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2" agemax="17" agemin="16" name="Kategorie B">
                  <RANKINGS>
                    <RANKING place="8" resultid="104" />
                    <RANKING place="4" resultid="265" />
                    <RANKING place="9" resultid="366" />
                    <RANKING place="2" resultid="637" />
                    <RANKING place="7" resultid="687" />
                    <RANKING place="6" resultid="723" />
                    <RANKING place="1" resultid="799" />
                    <RANKING place="3" resultid="926" />
                    <RANKING place="5" resultid="1084" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1" agemax="21" agemin="18" name="Junior:innen">
                  <RANKINGS>
                    <RANKING place="13" resultid="162" />
                    <RANKING place="12" resultid="189" />
                    <RANKING place="3" resultid="319" />
                    <RANKING place="2" resultid="432" />
                    <RANKING place="5" resultid="478" />
                    <RANKING place="1" resultid="680" />
                    <RANKING place="7" resultid="695" />
                    <RANKING place="14" resultid="713" />
                    <RANKING place="11" resultid="863" />
                    <RANKING place="9" resultid="1204" />
                    <RANKING place="8" resultid="1223" />
                    <RANKING place="10" resultid="1262" />
                    <RANKING place="6" resultid="1266" />
                    <RANKING place="4" resultid="1349" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="34" agemin="29" name="Master A">
                  <RANKINGS>
                    <RANKING place="1" resultid="969" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6" agemax="44" agemin="35" name="Master B">
                  <RANKINGS>
                    <RANKING place="1" resultid="70" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="7" agemax="54" agemin="45" name="Master C">
                  <RANKINGS>
                    <RANKING place="3" resultid="184" />
                    <RANKING place="5" resultid="542" />
                    <RANKING place="4" resultid="612" />
                    <RANKING place="9" resultid="646" />
                    <RANKING place="1" resultid="784" />
                    <RANKING place="7" resultid="803" />
                    <RANKING place="2" resultid="893" />
                    <RANKING place="6" resultid="1005" />
                    <RANKING place="8" resultid="1016" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8" agemax="64" agemin="55" name="Master D">
                  <RANKINGS>
                    <RANKING place="1" resultid="16" />
                    <RANKING place="3" resultid="58" />
                    <RANKING place="2" resultid="481" />
                    <RANKING place="4" resultid="830" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9" agemax="-1" agemin="65" name="Master E">
                  <RANKINGS>
                    <RANKING place="1" resultid="196" />
                    <RANKING place="2" resultid="1322" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10" agemax="-1" agemin="14" name="offene Wertung">
                  <RANKINGS>
                    <RANKING place="25" resultid="16" />
                    <RANKING place="54" resultid="58" />
                    <RANKING place="28" resultid="70" />
                    <RANKING place="41" resultid="104" />
                    <RANKING place="56" resultid="132" />
                    <RANKING place="40" resultid="139" />
                    <RANKING place="30" resultid="162" />
                    <RANKING place="39" resultid="184" />
                    <RANKING place="27" resultid="189" />
                    <RANKING place="53" resultid="196" />
                    <RANKING place="13" resultid="265" />
                    <RANKING place="10" resultid="319" />
                    <RANKING place="45" resultid="366" />
                    <RANKING place="58" resultid="402" />
                    <RANKING place="8" resultid="432" />
                    <RANKING place="35" resultid="453" />
                    <RANKING place="12" resultid="478" />
                    <RANKING place="50" resultid="481" />
                    <RANKING place="49" resultid="511" />
                    <RANKING place="43" resultid="526" />
                    <RANKING place="20" resultid="530" />
                    <RANKING place="46" resultid="542" />
                    <RANKING place="7" resultid="559" />
                    <RANKING place="44" resultid="603" />
                    <RANKING place="42" resultid="612" />
                    <RANKING place="4" resultid="637" />
                    <RANKING place="59" resultid="646" />
                    <RANKING place="6" resultid="680" />
                    <RANKING place="60" resultid="682" />
                    <RANKING place="36" resultid="687" />
                    <RANKING place="16" resultid="695" />
                    <RANKING place="61" resultid="697" />
                    <RANKING place="34" resultid="713" />
                    <RANKING place="18" resultid="719" />
                    <RANKING place="28" resultid="723" />
                    <RANKING place="31" resultid="784" />
                    <RANKING place="2" resultid="799" />
                    <RANKING place="51" resultid="803" />
                    <RANKING place="57" resultid="830" />
                    <RANKING place="55" resultid="852" />
                    <RANKING place="24" resultid="863" />
                    <RANKING place="22" resultid="890" />
                    <RANKING place="36" resultid="893" />
                    <RANKING place="32" resultid="919" />
                    <RANKING place="9" resultid="926" />
                    <RANKING place="3" resultid="949" />
                    <RANKING place="1" resultid="969" />
                    <RANKING place="47" resultid="1005" />
                    <RANKING place="52" resultid="1016" />
                    <RANKING place="26" resultid="1084" />
                    <RANKING place="47" resultid="1107" />
                    <RANKING place="14" resultid="1125" />
                    <RANKING place="38" resultid="1169" />
                    <RANKING place="33" resultid="1200" />
                    <RANKING place="19" resultid="1204" />
                    <RANKING place="17" resultid="1223" />
                    <RANKING place="21" resultid="1262" />
                    <RANKING place="15" resultid="1266" />
                    <RANKING place="62" resultid="1293" />
                    <RANKING place="63" resultid="1322" />
                    <RANKING place="11" resultid="1349" />
                    <RANKING place="23" resultid="1354" />
                    <RANKING place="5" resultid="1362" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11" agemax="-1" agemin="14" name="Internationale offene Wertung">
                  <RANKINGS>
                    <RANKING place="26" resultid="16" />
                    <RANKING place="56" resultid="58" />
                    <RANKING place="30" resultid="70" />
                    <RANKING place="43" resultid="104" />
                    <RANKING place="58" resultid="132" />
                    <RANKING place="42" resultid="139" />
                    <RANKING place="32" resultid="162" />
                    <RANKING place="41" resultid="184" />
                    <RANKING place="29" resultid="189" />
                    <RANKING place="55" resultid="196" />
                    <RANKING place="28" resultid="210" />
                    <RANKING place="13" resultid="265" />
                    <RANKING place="10" resultid="319" />
                    <RANKING place="47" resultid="366" />
                    <RANKING place="60" resultid="402" />
                    <RANKING place="8" resultid="432" />
                    <RANKING place="37" resultid="453" />
                    <RANKING place="12" resultid="478" />
                    <RANKING place="52" resultid="481" />
                    <RANKING place="51" resultid="511" />
                    <RANKING place="45" resultid="526" />
                    <RANKING place="20" resultid="530" />
                    <RANKING place="48" resultid="542" />
                    <RANKING place="7" resultid="559" />
                    <RANKING place="46" resultid="603" />
                    <RANKING place="44" resultid="612" />
                    <RANKING place="4" resultid="637" />
                    <RANKING place="61" resultid="646" />
                    <RANKING place="6" resultid="680" />
                    <RANKING place="62" resultid="682" />
                    <RANKING place="38" resultid="687" />
                    <RANKING place="16" resultid="695" />
                    <RANKING place="63" resultid="697" />
                    <RANKING place="36" resultid="713" />
                    <RANKING place="18" resultid="719" />
                    <RANKING place="30" resultid="723" />
                    <RANKING place="33" resultid="784" />
                    <RANKING place="2" resultid="799" />
                    <RANKING place="53" resultid="803" />
                    <RANKING place="59" resultid="830" />
                    <RANKING place="57" resultid="852" />
                    <RANKING place="25" resultid="863" />
                    <RANKING place="22" resultid="890" />
                    <RANKING place="38" resultid="893" />
                    <RANKING place="34" resultid="919" />
                    <RANKING place="9" resultid="926" />
                    <RANKING place="3" resultid="949" />
                    <RANKING place="1" resultid="969" />
                    <RANKING place="23" resultid="972" />
                    <RANKING place="49" resultid="1005" />
                    <RANKING place="54" resultid="1016" />
                    <RANKING place="27" resultid="1084" />
                    <RANKING place="49" resultid="1107" />
                    <RANKING place="14" resultid="1125" />
                    <RANKING place="40" resultid="1169" />
                    <RANKING place="35" resultid="1200" />
                    <RANKING place="19" resultid="1204" />
                    <RANKING place="17" resultid="1223" />
                    <RANKING place="21" resultid="1262" />
                    <RANKING place="15" resultid="1266" />
                    <RANKING place="64" resultid="1293" />
                    <RANKING place="65" resultid="1322" />
                    <RANKING place="11" resultid="1349" />
                    <RANKING place="24" resultid="1354" />
                    <RANKING place="5" resultid="1362" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="39" number="203" gender="F" round="TIM">
              <SWIMSTYLE stroke="BIFIN" relaycount="1" distance="50" />
              <FEE value="1000" currency="EUR" />
              <HEATS>
                <HEAT heatid="39001" number="1" />
                <HEAT heatid="39002" number="2" />
                <HEAT heatid="39003" number="3" />
                <HEAT heatid="39004" number="4" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="-1" agemin="12" name="offene Klasse">
                  <RANKINGS>
                    <RANKING place="5" resultid="81" />
                    <RANKING place="4" resultid="88" />
                    <RANKING place="16" resultid="217" />
                    <RANKING place="6" resultid="233" />
                    <RANKING place="22" resultid="396" />
                    <RANKING place="3" resultid="446" />
                    <RANKING place="9" resultid="458" />
                    <RANKING place="10" resultid="463" />
                    <RANKING place="11" resultid="521" />
                    <RANKING place="25" resultid="549" />
                    <RANKING place="8" resultid="582" />
                    <RANKING place="17" resultid="584" />
                    <RANKING place="13" resultid="656" />
                    <RANKING place="1" resultid="764" />
                    <RANKING place="21" resultid="835" />
                    <RANKING place="7" resultid="876" />
                    <RANKING place="20" resultid="895" />
                    <RANKING place="2" resultid="951" />
                    <RANKING place="26" resultid="995" />
                    <RANKING place="12" resultid="999" />
                    <RANKING place="14" resultid="1001" />
                    <RANKING place="15" resultid="1023" />
                    <RANKING place="19" resultid="1241" />
                    <RANKING place="24" resultid="1245" />
                    <RANKING place="23" resultid="1259" />
                    <RANKING place="18" resultid="1377" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="40" number="204" gender="M" round="TIM">
              <SWIMSTYLE stroke="BIFIN" relaycount="1" distance="50" />
              <FEE value="1000" currency="EUR" />
              <HEATS>
                <HEAT heatid="40001" number="1" />
                <HEAT heatid="40002" number="2" />
                <HEAT heatid="40003" number="3" />
                <HEAT heatid="40004" number="4" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemax="-1" agemin="12" name="offene Klasse">
                  <RANKINGS>
                    <RANKING place="17" resultid="18" />
                    <RANKING place="13" resultid="38" />
                    <RANKING place="2" resultid="166" />
                    <RANKING place="4" resultid="170" />
                    <RANKING place="14" resultid="186" />
                    <RANKING place="6" resultid="191" />
                    <RANKING place="5" resultid="212" />
                    <RANKING place="7" resultid="221" />
                    <RANKING place="15" resultid="483" />
                    <RANKING place="18" resultid="501" />
                    <RANKING place="19" resultid="513" />
                    <RANKING place="28" resultid="516" />
                    <RANKING place="27" resultid="544" />
                    <RANKING place="1" resultid="561" />
                    <RANKING place="20" resultid="683" />
                    <RANKING place="9" resultid="689" />
                    <RANKING place="12" resultid="714" />
                    <RANKING place="3" resultid="724" />
                    <RANKING place="25" resultid="741" />
                    <RANKING place="11" resultid="786" />
                    <RANKING place="21" resultid="805" />
                    <RANKING place="23" resultid="859" />
                    <RANKING place="10" resultid="973" />
                    <RANKING place="22" resultid="1003" />
                    <RANKING place="24" resultid="1007" />
                    <RANKING place="8" resultid="1013" />
                    <RANKING place="26" resultid="1018" />
                    <RANKING place="16" resultid="1027" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
          </EVENTS>
        </SESSION>
        <SESSION number="5" date="2023-05-14" daytime="15:37" officialmeeting="15:00" warmupfrom="14:30">
          <EVENTS>
            <EVENT eventid="41" number="117" gender="F" round="FIN">
              <SWIMSTYLE stroke="SURFACE" relaycount="1" distance="100" />
              <HEATS>
                <HEAT heatid="41000" number="0" />
                <HEAT heatid="41001" number="1" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="10" agemax="-1" agemin="12" name="offene Wertung">
                  <RANKINGS>
                    <RANKING place="2" resultid="1535" />
                    <RANKING place="7" resultid="1536" />
                    <RANKING place="1" resultid="1537" />
                    <RANKING place="4" resultid="1538" />
                    <RANKING place="3" resultid="1539" />
                    <RANKING place="6" resultid="1540" />
                    <RANKING place="5" resultid="1542" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11" agemax="-1" agemin="12" name="Internationale offene Wertung">
                  <RANKINGS>
                    <RANKING place="2" resultid="1535" />
                    <RANKING place="8" resultid="1536" />
                    <RANKING place="1" resultid="1537" />
                    <RANKING place="5" resultid="1538" />
                    <RANKING place="4" resultid="1539" />
                    <RANKING place="7" resultid="1540" />
                    <RANKING place="3" resultid="1541" />
                    <RANKING place="6" resultid="1542" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="42" number="118" gender="M" round="FIN">
              <SWIMSTYLE stroke="SURFACE" relaycount="1" distance="100" />
              <HEATS>
                <HEAT heatid="42001" number="1" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="10" agemax="-1" agemin="12" name="offene Wertung">
                  <RANKINGS>
                    <RANKING place="2" resultid="1543" />
                    <RANKING place="4" resultid="1544" />
                    <RANKING place="1" resultid="1545" />
                    <RANKING place="5" resultid="1546" />
                    <RANKING place="6" resultid="1547" />
                    <RANKING place="7" resultid="1548" />
                    <RANKING place="3" resultid="1549" />
                    <RANKING place="8" resultid="1550" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="43" number="319" gender="F" round="FIN">
              <SWIMSTYLE stroke="SURFACE" relaycount="1" distance="400" />
              <FEE value="650" currency="EUR" />
              <HEATS>
                <HEAT heatid="43001" number="1" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="4" agemax="13" agemin="12" name="Kategorie D" />
                <AGEGROUP agegroupid="3" agemax="15" agemin="14" name="Kategorie C" />
                <AGEGROUP agegroupid="2" agemax="17" agemin="16" name="Kategorie B">
                  <RANKINGS>
                    <RANKING place="2" resultid="428" />
                    <RANKING place="1" resultid="938" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1" agemax="21" agemin="18" name="Junior:innen">
                  <RANKINGS>
                    <RANKING place="3" resultid="770" />
                    <RANKING place="2" resultid="869" />
                    <RANKING place="1" resultid="1136" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="34" agemin="29" name="Master A" />
                <AGEGROUP agegroupid="6" agemax="44" agemin="35" name="Master B" />
                <AGEGROUP agegroupid="7" agemax="54" agemin="45" name="Master C" />
                <AGEGROUP agegroupid="8" agemax="64" agemin="55" name="Master D" />
                <AGEGROUP agegroupid="9" agemax="-1" agemin="65" name="Master E" />
                <AGEGROUP agegroupid="10" agemax="-1" agemin="12" name="offene Wertung">
                  <RANKINGS>
                    <RANKING place="4" resultid="428" />
                    <RANKING place="5" resultid="770" />
                    <RANKING place="3" resultid="869" />
                    <RANKING place="2" resultid="938" />
                    <RANKING place="1" resultid="1136" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11" agemax="-1" agemin="12" name="Internationale offene Wertung">
                  <RANKINGS>
                    <RANKING place="3" resultid="173" />
                    <RANKING place="5" resultid="428" />
                    <RANKING place="6" resultid="770" />
                    <RANKING place="4" resultid="869" />
                    <RANKING place="2" resultid="938" />
                    <RANKING place="1" resultid="1136" />
                    <RANKING place="7" resultid="1162" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="44" number="320" gender="M" round="FIN">
              <SWIMSTYLE stroke="SURFACE" relaycount="1" distance="400" />
              <FEE value="650" currency="EUR" />
              <HEATS>
                <HEAT heatid="44001" number="1" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="4" agemax="13" agemin="12" name="Kategorie D" />
                <AGEGROUP agegroupid="3" agemax="15" agemin="14" name="Kategorie C">
                  <RANKINGS>
                    <RANKING place="1" resultid="419" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2" agemax="17" agemin="16" name="Kategorie B">
                  <RANKINGS>
                    <RANKING place="1" resultid="925" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1" agemax="21" agemin="18" name="Junior:innen">
                  <RANKINGS>
                    <RANKING place="1" resultid="25" />
                    <RANKING place="3" resultid="391" />
                    <RANKING place="2" resultid="1265" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5" agemax="34" agemin="29" name="Master A" />
                <AGEGROUP agegroupid="6" agemax="44" agemin="35" name="Master B" />
                <AGEGROUP agegroupid="7" agemax="54" agemin="45" name="Master C" />
                <AGEGROUP agegroupid="8" agemax="64" agemin="55" name="Master D" />
                <AGEGROUP agegroupid="9" agemax="-1" agemin="65" name="Master E" />
                <AGEGROUP agegroupid="10" agemax="-1" agemin="12" name="offene Wertung">
                  <RANKINGS>
                    <RANKING place="3" resultid="25" />
                    <RANKING place="5" resultid="391" />
                    <RANKING place="6" resultid="419" />
                    <RANKING place="7" resultid="925" />
                    <RANKING place="1" resultid="933" />
                    <RANKING place="2" resultid="942" />
                    <RANKING place="4" resultid="1265" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11" agemax="-1" agemin="12" name="Internationale offene Wertung">
                  <RANKINGS>
                    <RANKING place="4" resultid="25" />
                    <RANKING place="6" resultid="391" />
                    <RANKING place="7" resultid="419" />
                    <RANKING place="8" resultid="925" />
                    <RANKING place="1" resultid="933" />
                    <RANKING place="3" resultid="942" />
                    <RANKING place="2" resultid="1174" />
                    <RANKING place="5" resultid="1265" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="45" number="123" gender="F" round="FIN">
              <SWIMSTYLE stroke="APNEA" relaycount="1" distance="50" />
              <HEATS>
                <HEAT heatid="45001" number="1" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="10" agemax="-1" agemin="12" name="offene Wertung">
                  <RANKINGS>
                    <RANKING place="1" resultid="1551" />
                    <RANKING place="3" resultid="1553" />
                    <RANKING place="5" resultid="1554" />
                    <RANKING place="4" resultid="1555" />
                    <RANKING place="6" resultid="1556" />
                    <RANKING place="2" resultid="1557" />
                    <RANKING place="7" resultid="1558" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11" agemax="-1" agemin="12" name="Internationale offene Wertung">
                  <RANKINGS>
                    <RANKING place="1" resultid="1551" />
                    <RANKING place="2" resultid="1552" />
                    <RANKING place="4" resultid="1553" />
                    <RANKING place="6" resultid="1554" />
                    <RANKING place="5" resultid="1555" />
                    <RANKING place="7" resultid="1556" />
                    <RANKING place="3" resultid="1557" />
                    <RANKING place="8" resultid="1558" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="46" number="124" gender="M" round="FIN">
              <SWIMSTYLE stroke="APNEA" relaycount="1" distance="50" />
              <HEATS>
                <HEAT heatid="46001" number="1" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="10" agemax="-1" agemin="12" name="offene Wertung">
                  <RANKINGS>
                    <RANKING place="2" resultid="1559" />
                    <RANKING place="1" resultid="1560" />
                    <RANKING place="3" resultid="1561" />
                    <RANKING place="4" resultid="1562" />
                    <RANKING place="5" resultid="1563" />
                    <RANKING place="6" resultid="1564" />
                    <RANKING place="7" resultid="1565" />
                    <RANKING place="8" resultid="1566" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="47" number="25" gender="X" round="TIM">
              <SWIMSTYLE stroke="SURFACE" relaycount="4" distance="100" />
              <FEE value="1000" currency="EUR" />
              <HEATS>
                <HEAT heatid="47001" number="1" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="5" agemax="-1" agemin="176" easy.ak="176" calculate="TOTAL" name="Master I" />
                <AGEGROUP agegroupid="6" agemax="-1" agemin="399" easy.ak="399" calculate="TOTAL" name="Master II">
                  <RANKINGS>
                    <RANKING place="1" resultid="2" />
                    <RANKING place="3" resultid="567" />
                    <RANKING place="4" resultid="820" />
                    <RANKING place="2" resultid="991" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="48" number="26" gender="F" round="TIM">
              <SWIMSTYLE stroke="SURFACE" relaycount="4" distance="100" />
              <FEE value="1000" currency="EUR" />
              <HEATS>
                <HEAT heatid="48001" number="1" />
                <HEAT heatid="48002" number="2" />
                <HEAT heatid="48003" number="3" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="4" agemax="13" agemin="12" name="Kategorie D">
                  <RANKINGS>
                    <RANKING place="1" resultid="816" />
                    <RANKING place="2" resultid="1337" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3" agemax="15" agemin="14" name="Kategorie C">
                  <RANKINGS>
                    <RANKING place="1" resultid="250" />
                    <RANKING place="3" resultid="409" />
                    <RANKING place="2" resultid="563" />
                    <RANKING place="4" resultid="1339" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2" agemax="17" agemin="16" name="Kategorie B">
                  <RANKINGS>
                    <RANKING place="5" resultid="359" />
                    <RANKING place="3" resultid="1184" />
                    <RANKING place="1" resultid="1330" />
                    <RANKING place="4" resultid="1333" />
                    <RANKING place="2" resultid="1376" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1" agemax="21" agemin="18" name="Junior:innen">
                  <RANKINGS>
                    <RANKING place="3" resultid="505" />
                    <RANKING place="2" resultid="817" />
                    <RANKING place="1" resultid="1112" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10" agemax="-1" agemin="12" name="offene Wertung">
                  <RANKINGS>
                    <RANKING place="10" resultid="134" />
                    <RANKING place="9" resultid="250" />
                    <RANKING place="13" resultid="359" />
                    <RANKING place="15" resultid="409" />
                    <RANKING place="7" resultid="505" />
                    <RANKING place="12" resultid="563" />
                    <RANKING place="14" resultid="816" />
                    <RANKING place="5" resultid="817" />
                    <RANKING place="2" resultid="908" />
                    <RANKING place="1" resultid="1112" />
                    <RANKING place="8" resultid="1184" />
                    <RANKING place="3" resultid="1330" />
                    <RANKING place="11" resultid="1333" />
                    <RANKING place="16" resultid="1337" />
                    <RANKING place="17" resultid="1339" />
                    <RANKING place="4" resultid="1376" />
                    <RANKING place="6" resultid="1383" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11" agemax="-1" agemin="12" name="Internationale offene Wertung">
                  <RANKINGS>
                    <RANKING place="12" resultid="134" />
                    <RANKING place="11" resultid="250" />
                    <RANKING place="15" resultid="359" />
                    <RANKING place="17" resultid="409" />
                    <RANKING place="9" resultid="505" />
                    <RANKING place="14" resultid="563" />
                    <RANKING place="16" resultid="816" />
                    <RANKING place="5" resultid="817" />
                    <RANKING place="2" resultid="908" />
                    <RANKING place="8" resultid="909" />
                    <RANKING place="1" resultid="1112" />
                    <RANKING place="7" resultid="1115" />
                    <RANKING place="10" resultid="1184" />
                    <RANKING place="3" resultid="1330" />
                    <RANKING place="13" resultid="1333" />
                    <RANKING place="18" resultid="1337" />
                    <RANKING place="19" resultid="1339" />
                    <RANKING place="4" resultid="1376" />
                    <RANKING place="6" resultid="1383" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="49" number="27" gender="M" round="TIM">
              <SWIMSTYLE stroke="SURFACE" relaycount="4" distance="100" />
              <FEE value="1000" currency="EUR" />
              <HEATS>
                <HEAT heatid="49001" number="1" />
                <HEAT heatid="49002" number="2" />
              </HEATS>
              <AGEGROUPS>
                <AGEGROUP agegroupid="4" agemax="13" agemin="12" name="Kategorie D">
                  <RANKINGS>
                    <RANKING place="1" resultid="565" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3" agemax="15" agemin="14" name="Kategorie C">
                  <RANKINGS>
                    <RANKING place="1" resultid="664" />
                    <RANKING place="2" resultid="1335" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2" agemax="17" agemin="16" name="Kategorie B">
                  <RANKINGS>
                    <RANKING place="1" resultid="89" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1" agemax="21" agemin="18" name="Junior:innen">
                  <RANKINGS>
                    <RANKING place="4" resultid="254" />
                    <RANKING place="2" resultid="405" />
                    <RANKING place="3" resultid="666" />
                    <RANKING place="1" resultid="1327" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10" agemax="-1" agemin="12" name="offene Wertung">
                  <RANKINGS>
                    <RANKING place="8" resultid="89" />
                    <RANKING place="6" resultid="254" />
                    <RANKING place="4" resultid="405" />
                    <RANKING place="10" resultid="565" />
                    <RANKING place="9" resultid="664" />
                    <RANKING place="5" resultid="666" />
                    <RANKING place="7" resultid="813" />
                    <RANKING place="1" resultid="905" />
                    <RANKING place="3" resultid="1110" />
                    <RANKING place="2" resultid="1327" />
                    <RANKING place="11" resultid="1335" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
            </EVENT>
          </EVENTS>
        </SESSION>
      </SESSIONS>
      <CLUBS>
        <CLUB name="1. Chemnitzer Tauchverein e.V." nation="GER" region="20" code="0">
          <ATHLETES>
            <ATHLETE athleteid="101" birthdate="2010-01-01" gender="F" lastname="Schwarzer" firstname="Angelina Sophie" license="0">
              <RESULTS>
                <RESULT resultid="360" eventid="1" swimtime="00:00:25.16" lane="6" heatid="1005" />
                <RESULT resultid="361" eventid="13" swimtime="00:00:57.50" lane="7" heatid="13002" />
                <RESULT resultid="362" eventid="17" swimtime="00:09:38.10" lane="1" heatid="17002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:03.27" />
                    <SPLIT distance="200" swimtime="00:02:15.02" />
                    <SPLIT distance="300" swimtime="00:03:30.23" />
                    <SPLIT distance="400" swimtime="00:04:46.62" />
                    <SPLIT distance="500" swimtime="00:06:02.36" />
                    <SPLIT distance="600" swimtime="00:07:17.54" />
                    <SPLIT distance="700" swimtime="00:08:31.17" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="363" eventid="31" swimtime="00:00:53.16" lane="4" heatid="31006" />
                <RESULT resultid="364" eventid="35" swimtime="00:00:24.62" lane="3" heatid="35002" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="102" birthdate="2006-01-01" gender="M" lastname="Lorenz" firstname="Emil" license="0">
              <RESULTS>
                <RESULT resultid="365" eventid="32" status="DNS" swimtime="00:00:00.00" lane="7" heatid="32010" />
                <RESULT resultid="366" eventid="38" swimtime="00:00:21.30" lane="6" heatid="38009" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="103" birthdate="2010-01-01" gender="F" lastname="Siegert" firstname="Emilia" license="0">
              <RESULTS>
                <RESULT resultid="367" eventid="1" status="DNS" swimtime="00:00:00.00" lane="6" heatid="1003" />
                <RESULT resultid="368" eventid="15" status="DNS" swimtime="00:00:00.00" lane="5" heatid="15002" />
                <RESULT resultid="369" eventid="31" status="DNS" swimtime="00:00:00.00" lane="4" heatid="31003" />
                <RESULT resultid="370" eventid="39" status="DNS" swimtime="00:00:00.00" lane="5" heatid="39001" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="104" birthdate="2011-01-01" gender="F" lastname="Nisch" firstname="Hanna Maria" license="0">
              <RESULTS>
                <RESULT resultid="371" eventid="1" swimtime="00:00:26.26" lane="2" heatid="1004" />
                <RESULT resultid="372" eventid="13" swimtime="00:01:03.67" lane="8" heatid="13002" />
                <RESULT resultid="373" eventid="17" swimtime="00:10:26.09" lane="4" heatid="17001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:11.42" />
                    <SPLIT distance="200" swimtime="00:02:31.55" />
                    <SPLIT distance="300" swimtime="00:03:54.19" />
                    <SPLIT distance="400" swimtime="00:05:15.56" />
                    <SPLIT distance="500" swimtime="00:06:36.61" />
                    <SPLIT distance="600" swimtime="00:07:58.73" />
                    <SPLIT distance="700" swimtime="00:09:17.52" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="374" eventid="31" status="DSQ" swimtime="00:00:58.64" lane="3" heatid="31004" comment="Falscher Start." />
                <RESULT resultid="375" eventid="35" swimtime="00:00:27.70" lane="4" heatid="35001" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="105" birthdate="2008-01-01" gender="F" lastname="Franke" firstname="Jenny" license="0">
              <RESULTS>
                <RESULT resultid="376" eventid="1" swimtime="00:00:21.92" lane="3" heatid="1010" />
                <RESULT resultid="377" eventid="13" swimtime="00:00:53.02" lane="5" heatid="13003" />
                <RESULT resultid="378" eventid="17" swimtime="00:09:05.62" lane="6" heatid="17002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:58.34" />
                    <SPLIT distance="200" swimtime="00:02:05.02" />
                    <SPLIT distance="300" swimtime="00:03:14.48" />
                    <SPLIT distance="400" swimtime="00:04:25.50" />
                    <SPLIT distance="500" swimtime="00:05:36.53" />
                    <SPLIT distance="600" swimtime="00:06:48.36" />
                    <SPLIT distance="700" swimtime="00:07:59.15" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="379" eventid="31" swimtime="00:00:48.33" lane="3" heatid="31011" />
                <RESULT resultid="380" eventid="37" swimtime="00:00:19.76" lane="8" heatid="37004" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="106" birthdate="2007-01-01" gender="F" lastname="Ullrich" firstname="Johanna Hermine" license="0">
              <RESULTS>
                <RESULT resultid="381" eventid="3" swimtime="00:16:44.04" lane="6" heatid="3001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:56.49" />
                    <SPLIT distance="200" swimtime="00:02:01.53" />
                    <SPLIT distance="300" swimtime="00:03:09.69" />
                    <SPLIT distance="400" swimtime="00:04:18.29" />
                    <SPLIT distance="500" swimtime="00:05:26.46" />
                    <SPLIT distance="600" swimtime="00:06:36.62" />
                    <SPLIT distance="700" swimtime="00:07:45.88" />
                    <SPLIT distance="800" swimtime="00:08:53.96" />
                    <SPLIT distance="900" swimtime="00:10:02.83" />
                    <SPLIT distance="1000" swimtime="00:11:10.96" />
                    <SPLIT distance="1100" swimtime="00:12:20.30" />
                    <SPLIT distance="1200" swimtime="00:13:29.96" />
                    <SPLIT distance="1300" swimtime="00:14:38.30" />
                    <SPLIT distance="1400" swimtime="00:15:44.72" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="382" eventid="13" swimtime="00:00:53.16" lane="3" heatid="13003" />
                <RESULT resultid="383" eventid="17" swimtime="00:08:43.57" lane="4" heatid="17003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:55.37" />
                    <SPLIT distance="200" swimtime="00:02:02.49" />
                    <SPLIT distance="300" swimtime="00:03:09.57" />
                    <SPLIT distance="400" swimtime="00:04:18.55" />
                    <SPLIT distance="500" swimtime="00:05:27.44" />
                    <SPLIT distance="600" swimtime="00:06:36.38" />
                    <SPLIT distance="700" swimtime="00:07:43.31" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="384" eventid="33" swimtime="00:04:11.94" lane="8" heatid="33005">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:57.41" />
                    <SPLIT distance="200" swimtime="00:02:03.72" />
                    <SPLIT distance="300" swimtime="00:03:10.82" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="385" eventid="37" swimtime="00:00:22.98" lane="8" heatid="37002" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="107" birthdate="2005-01-01" gender="M" lastname="Porges" firstname="Marcel" license="0">
              <RESULTS>
                <RESULT resultid="386" eventid="2" swimtime="00:00:17.20" lane="5" heatid="2010" />
                <RESULT resultid="1416" eventid="8" swimtime="00:00:17.68" lane="2" heatid="8001" />
                <RESULT resultid="387" eventid="16" swimtime="00:01:31.83" lane="3" heatid="16007">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:44.28" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1522" eventid="24" status="WDR" swimtime="00:00:00.00" lane="0" heatid="24000" />
                <RESULT resultid="388" eventid="26" swimtime="00:07:11.49" lane="3" heatid="26001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:47.83" />
                    <SPLIT distance="200" swimtime="00:01:41.54" />
                    <SPLIT distance="300" swimtime="00:02:37.52" />
                    <SPLIT distance="400" swimtime="00:03:33.67" />
                    <SPLIT distance="500" swimtime="00:04:29.69" />
                    <SPLIT distance="600" swimtime="00:05:26.22" />
                    <SPLIT distance="700" swimtime="00:06:20.73" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="389" eventid="28" swimtime="00:03:11.34" lane="8" heatid="28001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:43.90" />
                    <SPLIT distance="200" swimtime="00:01:32.87" />
                    <SPLIT distance="300" swimtime="00:02:23.56" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="390" eventid="32" swimtime="00:00:40.01" lane="3" heatid="32012" />
                <RESULT resultid="1548" eventid="42" swimtime="00:00:40.37" lane="7" heatid="42001" />
                <RESULT resultid="391" eventid="44" swimtime="00:03:31.80" lane="7" heatid="44001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:48.41" />
                    <SPLIT distance="200" swimtime="00:01:40.91" />
                    <SPLIT distance="300" swimtime="00:02:36.52" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="108" birthdate="2010-01-01" gender="F" lastname="Bluhm" firstname="Suna" license="0">
              <RESULTS>
                <RESULT resultid="392" eventid="1" swimtime="00:00:28.56" lane="2" heatid="1002" />
                <RESULT resultid="395" eventid="5" swimtime="00:01:14.52" lane="1" heatid="5002" />
                <RESULT resultid="393" eventid="15" status="DSQ" swimtime="00:02:33.51" lane="4" heatid="15002" comment="Falscher Start.">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:14.64" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="394" eventid="31" swimtime="00:01:03.14" lane="1" heatid="31003" />
                <RESULT resultid="396" eventid="39" swimtime="00:00:31.26" lane="1" heatid="39001" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="109" birthdate="2009-01-01" gender="M" lastname="Hans" firstname="Yannick" license="0">
              <RESULTS>
                <RESULT resultid="397" eventid="2" swimtime="00:00:24.56" lane="8" heatid="2005" />
                <RESULT resultid="403" eventid="6" status="DSQ" swimtime="00:01:01.43" lane="2" heatid="6003" comment="Falscher Stil." />
                <RESULT resultid="398" eventid="16" swimtime="00:01:58.76" lane="4" heatid="16004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:56.69" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="399" eventid="18" swimtime="00:09:24.12" lane="8" heatid="18002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:02.92" />
                    <SPLIT distance="200" swimtime="00:02:14.59" />
                    <SPLIT distance="300" swimtime="00:03:26.72" />
                    <SPLIT distance="400" swimtime="00:04:39.40" />
                    <SPLIT distance="500" swimtime="00:05:53.67" />
                    <SPLIT distance="600" swimtime="00:07:08.46" />
                    <SPLIT distance="700" swimtime="00:08:22.00" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="400" eventid="32" swimtime="00:00:53.67" lane="7" heatid="32005" />
                <RESULT resultid="401" eventid="34" swimtime="00:04:17.71" lane="1" heatid="34005">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:57.96" />
                    <SPLIT distance="200" swimtime="00:02:06.41" />
                    <SPLIT distance="300" swimtime="00:03:16.10" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="402" eventid="38" swimtime="00:00:24.16" lane="7" heatid="38003" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY number="1" gender="F" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="358" eventid="11" swimtime="00:08:16.14" lane="5" heatid="11001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:59.47" />
                    <SPLIT distance="200" swimtime="00:02:06.53" />
                    <SPLIT distance="300" swimtime="00:03:01.86" />
                    <SPLIT distance="400" swimtime="00:04:02.96" />
                    <SPLIT distance="500" swimtime="00:05:10.28" />
                    <SPLIT distance="600" swimtime="00:06:24.16" />
                    <SPLIT distance="700" swimtime="00:07:16.46" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="101" number="1" />
                    <RELAYPOSITION athleteid="106" number="2" />
                    <RELAYPOSITION athleteid="104" number="3" />
                    <RELAYPOSITION athleteid="105" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="2" gender="F" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="359" eventid="48" swimtime="00:03:39.64" lane="1" heatid="48002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:53.05" />
                    <SPLIT distance="200" swimtime="00:01:49.74" />
                    <SPLIT distance="300" swimtime="00:02:51.52" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="106" number="1" />
                    <RELAYPOSITION athleteid="101" number="2" />
                    <RELAYPOSITION athleteid="104" number="3" />
                    <RELAYPOSITION athleteid="105" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB name="Aquanauten Karlsruhe-Durlach e.V." nation="GER" region="33" code="0">
          <ATHLETES>
            <ATHLETE athleteid="10" birthdate="2007-01-01" gender="F" lastname="Kirchner" firstname="Nia" license="0">
              <RESULTS>
                <RESULT resultid="50" eventid="1" swimtime="00:00:22.95" lane="5" heatid="1007" />
                <RESULT resultid="51" eventid="3" swimtime="00:16:39.65" lane="1" heatid="3002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:58.91" />
                    <SPLIT distance="200" swimtime="00:02:03.62" />
                    <SPLIT distance="300" swimtime="00:03:11.46" />
                    <SPLIT distance="400" swimtime="00:04:17.14" />
                    <SPLIT distance="500" swimtime="00:05:25.24" />
                    <SPLIT distance="600" swimtime="00:06:33.23" />
                    <SPLIT distance="700" swimtime="00:07:42.16" />
                    <SPLIT distance="800" swimtime="00:08:50.65" />
                    <SPLIT distance="900" swimtime="00:10:01.24" />
                    <SPLIT distance="1000" swimtime="00:11:11.29" />
                    <SPLIT distance="1100" swimtime="00:12:19.38" />
                    <SPLIT distance="1200" swimtime="00:13:29.58" />
                    <SPLIT distance="1300" swimtime="00:14:38.52" />
                    <SPLIT distance="1400" swimtime="00:15:42.40" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="52" eventid="13" swimtime="00:00:49.96" lane="7" heatid="13004" />
                <RESULT resultid="53" eventid="17" swimtime="00:08:18.96" lane="5" heatid="17004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:56.88" />
                    <SPLIT distance="200" swimtime="00:02:01.83" />
                    <SPLIT distance="300" swimtime="00:03:07.82" />
                    <SPLIT distance="400" swimtime="00:04:13.22" />
                    <SPLIT distance="500" swimtime="00:05:16.36" />
                    <SPLIT distance="600" swimtime="00:06:21.33" />
                    <SPLIT distance="700" swimtime="00:07:24.42" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="Berliner TSC e.V." nation="GER" region="21" code="304088">
          <ATHLETES>
            <ATHLETE athleteid="115" birthdate="2009-01-01" gender="F" lastname="Grabner" firstname="Anabel" license="0">
              <RESULTS>
                <RESULT resultid="411" eventid="1" swimtime="00:00:25.91" lane="3" heatid="1003" />
                <RESULT resultid="412" eventid="15" swimtime="00:02:04.87" lane="6" heatid="15004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:00.79" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="413" eventid="31" swimtime="00:00:57.96" lane="6" heatid="31004" />
                <RESULT resultid="414" eventid="33" swimtime="00:04:35.15" lane="5" heatid="33002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:06.17" />
                    <SPLIT distance="200" swimtime="00:02:18.27" />
                    <SPLIT distance="300" swimtime="00:03:31.07" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="116" birthdate="2008-01-01" gender="M" lastname="Welke" firstname="Anton" license="0">
              <RESULTS>
                <RESULT resultid="415" eventid="2" swimtime="00:00:20.19" lane="8" heatid="2011" />
                <RESULT resultid="416" eventid="16" swimtime="00:01:38.69" lane="6" heatid="16006">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:46.13" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="417" eventid="26" swimtime="00:07:26.98" lane="7" heatid="26001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:49.93" />
                    <SPLIT distance="200" swimtime="00:01:46.92" />
                    <SPLIT distance="300" swimtime="00:02:43.88" />
                    <SPLIT distance="400" swimtime="00:03:41.46" />
                    <SPLIT distance="500" swimtime="00:04:38.43" />
                    <SPLIT distance="600" swimtime="00:05:35.70" />
                    <SPLIT distance="700" swimtime="00:06:32.63" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="418" eventid="32" status="DSQ" swimtime="00:00:43.73" lane="8" heatid="32011" comment="Falscher Start." />
                <RESULT resultid="419" eventid="44" swimtime="00:03:37.61" lane="8" heatid="44001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:49.96" />
                    <SPLIT distance="200" swimtime="00:01:45.35" />
                    <SPLIT distance="300" swimtime="00:02:42.22" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="117" birthdate="2011-01-01" gender="F" lastname="Stobbe" firstname="Bella" license="123">
              <RESULTS>
                <RESULT resultid="420" eventid="3" swimtime="00:19:25.02" lane="2" heatid="3001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:09.26" />
                    <SPLIT distance="200" swimtime="00:02:26.78" />
                    <SPLIT distance="300" swimtime="00:03:45.05" />
                    <SPLIT distance="400" swimtime="00:05:03.66" />
                    <SPLIT distance="500" swimtime="00:06:22.51" />
                    <SPLIT distance="600" swimtime="00:07:41.91" />
                    <SPLIT distance="700" swimtime="00:09:01.84" />
                    <SPLIT distance="800" swimtime="00:10:21.95" />
                    <SPLIT distance="900" swimtime="00:11:40.57" />
                    <SPLIT distance="1000" swimtime="00:12:59.99" />
                    <SPLIT distance="1100" swimtime="00:14:19.58" />
                    <SPLIT distance="1200" swimtime="00:15:38.22" />
                    <SPLIT distance="1300" swimtime="00:16:57.05" />
                    <SPLIT distance="1400" swimtime="00:18:11.75" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="421" eventid="17" swimtime="00:09:08.38" lane="6" heatid="17003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:02.76" />
                    <SPLIT distance="200" swimtime="00:02:12.09" />
                    <SPLIT distance="300" swimtime="00:03:21.83" />
                    <SPLIT distance="400" swimtime="00:04:31.96" />
                    <SPLIT distance="500" swimtime="00:05:43.82" />
                    <SPLIT distance="600" swimtime="00:06:54.21" />
                    <SPLIT distance="700" swimtime="00:08:02.50" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="422" eventid="31" swimtime="00:00:58.86" lane="7" heatid="31006" />
                <RESULT resultid="423" eventid="33" swimtime="00:04:26.03" lane="5" heatid="33003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:02.43" />
                    <SPLIT distance="200" swimtime="00:02:11.48" />
                    <SPLIT distance="300" swimtime="00:03:21.15" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="118" birthdate="2007-01-01" gender="F" lastname="Eggert" firstname="Emilia" license="0">
              <RESULTS>
                <RESULT resultid="424" eventid="1" swimtime="00:00:20.40" lane="1" heatid="1015" />
                <RESULT resultid="425" eventid="15" swimtime="00:01:39.33" lane="3" heatid="15010">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:47.48" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1512" eventid="23" status="WDR" swimtime="00:00:00.00" lane="0" heatid="23000" />
                <RESULT resultid="426" eventid="27" swimtime="00:03:38.83" lane="2" heatid="27001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:50.95" />
                    <SPLIT distance="200" swimtime="00:01:46.33" />
                    <SPLIT distance="300" swimtime="00:02:43.58" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="427" eventid="31" swimtime="00:00:45.18" lane="6" heatid="31017" />
                <RESULT resultid="429" eventid="37" swimtime="00:00:19.02" lane="6" heatid="37007" />
                <RESULT resultid="1533" eventid="41" status="WDR" swimtime="00:00:00.00" lane="0" heatid="41000" />
                <RESULT resultid="428" eventid="43" swimtime="00:03:39.67" lane="2" heatid="43001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:49.89" />
                    <SPLIT distance="200" swimtime="00:01:45.56" />
                    <SPLIT distance="300" swimtime="00:02:43.45" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="119" birthdate="2005-01-01" gender="M" lastname="Bandlow" firstname="Jan" license="0">
              <RESULTS>
                <RESULT resultid="430" eventid="2" swimtime="00:00:19.45" lane="8" heatid="2009" />
                <RESULT resultid="431" eventid="32" swimtime="00:00:43.76" lane="2" heatid="32009" />
                <RESULT resultid="432" eventid="38" swimtime="00:00:17.00" lane="2" heatid="38009" />
                <RESULT resultid="1566" eventid="46" swimtime="00:00:16.95" lane="8" heatid="46001" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="120" birthdate="2007-01-01" gender="F" lastname="Beske" firstname="Lena" license="0">
              <RESULTS>
                <RESULT resultid="433" eventid="1" swimtime="00:00:23.76" lane="8" heatid="1011" />
                <RESULT resultid="434" eventid="13" swimtime="00:00:53.12" lane="4" heatid="13003" />
                <RESULT resultid="435" eventid="31" swimtime="00:00:52.96" lane="2" heatid="31010" />
                <RESULT resultid="436" eventid="37" swimtime="00:00:21.06" lane="8" heatid="37005" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="121" birthdate="2009-01-01" gender="F" lastname="Herzog" firstname="Matilda" license="123">
              <RESULTS>
                <RESULT resultid="437" eventid="1" swimtime="00:00:24.06" lane="2" heatid="1008" />
                <RESULT resultid="438" eventid="15" swimtime="00:01:59.50" lane="1" heatid="15007">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:57.96" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="439" eventid="31" swimtime="00:00:53.71" lane="4" heatid="31009" />
                <RESULT resultid="440" eventid="33" swimtime="00:04:15.02" lane="6" heatid="33004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:00.31" />
                    <SPLIT distance="200" swimtime="00:02:08.51" />
                    <SPLIT distance="300" swimtime="00:03:14.65" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="122" birthdate="2007-01-01" gender="F" lastname="Manthey" firstname="Maxime" license="123">
              <RESULTS>
                <RESULT resultid="441" eventid="1" swimtime="00:00:20.05" lane="6" heatid="1014" />
                <RESULT resultid="442" eventid="13" swimtime="00:00:41.60" lane="3" heatid="13007" />
                <RESULT resultid="443" eventid="15" swimtime="00:01:44.87" lane="6" heatid="15012">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:49.29" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1499" eventid="21" swimtime="00:00:42.11" lane="1" heatid="21001" />
                <RESULT resultid="444" eventid="31" swimtime="00:00:46.01" lane="2" heatid="31016" />
                <RESULT resultid="445" eventid="37" swimtime="00:00:17.92" lane="5" heatid="37008" />
                <RESULT resultid="446" eventid="39" swimtime="00:00:24.04" lane="3" heatid="39004" />
                <RESULT resultid="1554" eventid="45" swimtime="00:00:18.09" lane="6" heatid="45001" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="123" birthdate="2009-10-17" gender="F" lastname="Chelius" firstname="Nahla" license="123">
              <RESULTS>
                <RESULT resultid="447" eventid="31" swimtime="00:00:59.74" lane="5" heatid="31004" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="124" birthdate="2009-01-01" gender="M" lastname="Martiny" firstname="Peter" license="0">
              <RESULTS>
                <RESULT resultid="448" eventid="4" swimtime="00:16:01.77" lane="6" heatid="4001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:52.41" />
                    <SPLIT distance="200" swimtime="00:01:55.45" />
                    <SPLIT distance="300" swimtime="00:03:01.73" />
                    <SPLIT distance="400" swimtime="00:04:06.78" />
                    <SPLIT distance="500" swimtime="00:05:12.32" />
                    <SPLIT distance="600" swimtime="00:06:18.73" />
                    <SPLIT distance="700" swimtime="00:07:23.29" />
                    <SPLIT distance="800" swimtime="00:08:29.83" />
                    <SPLIT distance="900" swimtime="00:09:35.09" />
                    <SPLIT distance="1000" swimtime="00:10:40.46" />
                    <SPLIT distance="1100" swimtime="00:11:45.84" />
                    <SPLIT distance="1200" swimtime="00:12:51.51" />
                    <SPLIT distance="1300" swimtime="00:13:58.33" />
                    <SPLIT distance="1400" swimtime="00:15:02.07" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="449" eventid="16" swimtime="00:01:49.13" lane="1" heatid="16003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:50.07" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="450" eventid="26" swimtime="00:08:06.27" lane="8" heatid="26001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:52.91" />
                    <SPLIT distance="200" swimtime="00:01:53.79" />
                    <SPLIT distance="300" swimtime="00:02:57.01" />
                    <SPLIT distance="400" swimtime="00:04:00.56" />
                    <SPLIT distance="500" swimtime="00:05:04.10" />
                    <SPLIT distance="600" swimtime="00:06:06.72" />
                    <SPLIT distance="700" swimtime="00:07:08.36" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="451" eventid="32" swimtime="00:00:48.01" lane="4" heatid="32007" />
                <RESULT resultid="452" eventid="34" swimtime="00:03:56.92" lane="7" heatid="34006">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:53.03" />
                    <SPLIT distance="200" swimtime="00:01:56.08" />
                    <SPLIT distance="300" swimtime="00:02:59.20" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="453" eventid="38" swimtime="00:00:20.18" lane="5" heatid="38004" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="125" birthdate="2003-01-01" gender="F" lastname="Fränzel" firstname="Samirah" license="123">
              <RESULTS>
                <RESULT resultid="454" eventid="1" swimtime="00:00:22.04" lane="1" heatid="1009" />
                <RESULT resultid="457" eventid="5" swimtime="00:00:59.58" lane="3" heatid="5003" />
                <RESULT resultid="455" eventid="31" swimtime="00:00:50.94" lane="8" heatid="31010" />
                <RESULT resultid="456" eventid="37" swimtime="00:00:21.52" lane="5" heatid="37002" />
                <RESULT resultid="458" eventid="39" swimtime="00:00:26.44" lane="6" heatid="39003" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="126" birthdate="2009-05-26" gender="F" lastname="Ivanova" firstname="Taisiia" license="123">
              <RESULTS>
                <RESULT resultid="459" eventid="1" swimtime="00:00:25.05" lane="2" heatid="1007" />
                <RESULT resultid="462" eventid="5" swimtime="00:01:01.79" lane="1" heatid="5003" />
                <RESULT resultid="460" eventid="15" swimtime="00:02:07.60" lane="5" heatid="15004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:01.55" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="461" eventid="31" swimtime="00:00:57.33" lane="2" heatid="31007" />
                <RESULT resultid="463" eventid="39" swimtime="00:00:27.24" lane="5" heatid="39002" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="127" birthdate="2008-01-01" gender="F" lastname="Bublitz" firstname="Tessa" license="123">
              <RESULTS>
                <RESULT resultid="464" eventid="1" swimtime="00:00:21.42" lane="7" heatid="1014" />
                <RESULT resultid="465" eventid="15" swimtime="00:01:45.92" lane="7" heatid="15012">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:49.99" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="466" eventid="25" swimtime="00:07:51.29" lane="2" heatid="25001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:53.82" />
                    <SPLIT distance="200" swimtime="00:01:53.19" />
                    <SPLIT distance="300" swimtime="00:02:54.56" />
                    <SPLIT distance="400" swimtime="00:03:55.27" />
                    <SPLIT distance="500" swimtime="00:04:56.32" />
                    <SPLIT distance="600" swimtime="00:05:57.39" />
                    <SPLIT distance="700" swimtime="00:06:56.43" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="467" eventid="31" swimtime="00:00:47.73" lane="7" heatid="31016" />
                <RESULT resultid="468" eventid="33" swimtime="00:03:46.31" lane="4" heatid="33007">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:51.48" />
                    <SPLIT distance="200" swimtime="00:01:50.83" />
                    <SPLIT distance="300" swimtime="00:02:50.60" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="469" eventid="37" swimtime="00:00:20.15" lane="8" heatid="37006" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="129" birthdate="2004-01-01" gender="M" lastname="Beske" firstname="Tom" license="0">
              <RESULTS>
                <RESULT resultid="474" eventid="2" swimtime="00:00:18.63" lane="6" heatid="2011" />
                <RESULT resultid="475" eventid="14" swimtime="00:00:37.92" lane="5" heatid="14005" />
                <RESULT resultid="1508" eventid="22" swimtime="00:00:37.92" lane="2" heatid="22001" />
                <RESULT resultid="476" eventid="28" swimtime="00:03:10.03" lane="4" heatid="28001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:42.94" />
                    <SPLIT distance="200" swimtime="00:01:30.29" />
                    <SPLIT distance="300" swimtime="00:02:21.56" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="477" eventid="32" swimtime="00:00:39.49" lane="3" heatid="32010" />
                <RESULT resultid="478" eventid="38" swimtime="00:00:17.20" lane="2" heatid="38008" />
                <RESULT resultid="1547" eventid="42" swimtime="00:00:39.10" lane="2" heatid="42001" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY number="1" gender="M" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="404" eventid="12" swimtime="00:06:48.70" lane="6" heatid="12002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:46.28" />
                    <SPLIT distance="200" swimtime="00:01:40.63" />
                    <SPLIT distance="300" swimtime="00:02:26.12" />
                    <SPLIT distance="400" swimtime="00:03:25.36" />
                    <SPLIT distance="500" swimtime="00:04:15.90" />
                    <SPLIT distance="600" swimtime="00:05:05.61" />
                    <SPLIT distance="700" swimtime="00:05:58.53" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="116" number="1" />
                    <RELAYPOSITION athleteid="119" number="2" />
                    <RELAYPOSITION athleteid="124" number="3" />
                    <RELAYPOSITION athleteid="129" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT resultid="405" eventid="49" swimtime="00:02:54.68" lane="6" heatid="49002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:40.10" />
                    <SPLIT distance="200" swimtime="00:01:23.23" />
                    <SPLIT distance="300" swimtime="00:02:11.21" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="129" number="1" />
                    <RELAYPOSITION athleteid="119" number="2" />
                    <RELAYPOSITION athleteid="124" number="3" />
                    <RELAYPOSITION athleteid="116" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" gender="F" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="406" eventid="11" swimtime="00:07:08.60" lane="2" heatid="11003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:47.38" />
                    <SPLIT distance="200" swimtime="00:01:39.22" />
                    <SPLIT distance="300" swimtime="00:02:30.01" />
                    <SPLIT distance="400" swimtime="00:03:26.32" />
                    <SPLIT distance="500" swimtime="00:04:21.72" />
                    <SPLIT distance="600" swimtime="00:05:24.31" />
                    <SPLIT distance="700" swimtime="00:06:12.52" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="118" number="1" />
                    <RELAYPOSITION athleteid="127" number="2" />
                    <RELAYPOSITION athleteid="121" number="3" />
                    <RELAYPOSITION athleteid="122" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" gender="X" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="408" eventid="30" swimtime="00:01:16.32" lane="6" heatid="30004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:38.38" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="122" number="1" />
                    <RELAYPOSITION athleteid="119" number="2" />
                    <RELAYPOSITION athleteid="118" number="3" />
                    <RELAYPOSITION athleteid="129" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="2" gender="F" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="409" eventid="48" swimtime="00:03:48.74" lane="4" heatid="48001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:58.45" />
                    <SPLIT distance="200" swimtime="00:01:56.76" />
                    <SPLIT distance="300" swimtime="00:02:55.04" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="117" number="1" />
                    <RELAYPOSITION athleteid="115" number="2" />
                    <RELAYPOSITION athleteid="123" number="3" />
                    <RELAYPOSITION athleteid="121" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="2" gender="X" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="410" eventid="30" swimtime="00:01:25.20" lane="2" heatid="30003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:42.29" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="124" number="1" />
                    <RELAYPOSITION athleteid="127" number="2" />
                    <RELAYPOSITION athleteid="121" number="3" />
                    <RELAYPOSITION athleteid="116" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" gender="F" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="1376" eventid="48" swimtime="00:03:09.98" lane="7" heatid="48003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:45.87" />
                    <SPLIT distance="200" swimtime="00:01:33.29" />
                    <SPLIT distance="300" swimtime="00:02:25.95" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="122" number="1" />
                    <RELAYPOSITION athleteid="127" number="2" />
                    <RELAYPOSITION athleteid="120" number="3" />
                    <RELAYPOSITION athleteid="118" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB name="Binger Tauchsportclub e.V." nation="GER" region="29" code="0">
          <ATHLETES>
            <ATHLETE athleteid="38" birthdate="2010-01-01" gender="M" lastname="Funke" firstname="Florian" license="0">
              <RESULTS>
                <RESULT resultid="92" eventid="2" swimtime="00:00:26.16" lane="1" heatid="2004" />
                <RESULT resultid="93" eventid="4" swimtime="00:21:00.74" lane="3" heatid="4001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:15.97" />
                    <SPLIT distance="200" swimtime="00:02:38.59" />
                    <SPLIT distance="300" swimtime="00:03:59.70" />
                    <SPLIT distance="400" swimtime="00:05:23.35" />
                    <SPLIT distance="500" swimtime="00:06:48.36" />
                    <SPLIT distance="600" swimtime="00:08:13.91" />
                    <SPLIT distance="700" swimtime="00:09:38.92" />
                    <SPLIT distance="800" swimtime="00:11:05.25" />
                    <SPLIT distance="900" swimtime="00:12:29.75" />
                    <SPLIT distance="1000" swimtime="00:13:53.82" />
                    <SPLIT distance="1100" swimtime="00:15:21.46" />
                    <SPLIT distance="1200" swimtime="00:16:51.18" />
                    <SPLIT distance="1300" swimtime="00:18:22.92" />
                    <SPLIT distance="1400" swimtime="00:19:46.51" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="94" eventid="16" swimtime="00:02:13.86" lane="8" heatid="16004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:03.62" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="95" eventid="18" swimtime="00:09:47.40" lane="2" heatid="18002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:11.23" />
                    <SPLIT distance="200" swimtime="00:02:28.46" />
                    <SPLIT distance="300" swimtime="00:03:44.21" />
                    <SPLIT distance="400" swimtime="00:04:57.72" />
                    <SPLIT distance="500" swimtime="00:06:10.12" />
                    <SPLIT distance="600" swimtime="00:07:23.58" />
                    <SPLIT distance="700" swimtime="00:08:35.79" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="96" eventid="32" swimtime="00:00:58.07" lane="6" heatid="32003" />
                <RESULT resultid="97" eventid="34" swimtime="00:04:36.01" lane="4" heatid="34003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:06.36" />
                    <SPLIT distance="200" swimtime="00:02:16.74" />
                    <SPLIT distance="300" swimtime="00:03:27.07" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="39" birthdate="2006-01-01" gender="M" lastname="Blaszczyk" firstname="Jan" license="0">
              <RESULTS>
                <RESULT resultid="98" eventid="2" status="DNS" swimtime="00:00:00.00" lane="4" heatid="2007" />
                <RESULT resultid="105" eventid="6" swimtime="00:00:57.96" lane="6" heatid="6002" />
                <RESULT resultid="99" eventid="14" swimtime="00:00:52.72" lane="8" heatid="14003" />
                <RESULT resultid="100" eventid="16" swimtime="00:01:54.78" lane="2" heatid="16005">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:55.56" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="101" eventid="18" swimtime="00:08:47.09" lane="6" heatid="18003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:00.47" />
                    <SPLIT distance="200" swimtime="00:02:05.94" />
                    <SPLIT distance="300" swimtime="00:03:12.33" />
                    <SPLIT distance="400" swimtime="00:04:19.34" />
                    <SPLIT distance="500" swimtime="00:05:26.23" />
                    <SPLIT distance="600" swimtime="00:06:32.67" />
                    <SPLIT distance="700" swimtime="00:07:35.09" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="102" eventid="32" swimtime="00:00:49.48" lane="7" heatid="32007" />
                <RESULT resultid="103" eventid="34" swimtime="00:04:07.09" lane="7" heatid="34005">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:55.72" />
                    <SPLIT distance="200" swimtime="00:01:58.44" />
                    <SPLIT distance="300" swimtime="00:03:03.53" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="104" eventid="38" swimtime="00:00:20.84" lane="4" heatid="38004" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="40" birthdate="2004-01-01" gender="F" lastname="Walter" firstname="Julia" license="0">
              <RESULTS>
                <RESULT resultid="106" eventid="1" swimtime="00:00:22.95" lane="8" heatid="1009" />
                <RESULT resultid="107" eventid="9" swimtime="00:16:38.94" lane="8" heatid="9001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:56.08" />
                    <SPLIT distance="200" swimtime="00:01:58.95" />
                    <SPLIT distance="300" swimtime="00:03:04.42" />
                    <SPLIT distance="400" swimtime="00:04:11.28" />
                    <SPLIT distance="500" swimtime="00:05:17.87" />
                    <SPLIT distance="600" swimtime="00:06:25.90" />
                    <SPLIT distance="700" swimtime="00:07:34.73" />
                    <SPLIT distance="800" swimtime="00:08:43.43" />
                    <SPLIT distance="900" swimtime="00:09:52.29" />
                    <SPLIT distance="1000" swimtime="00:11:01.84" />
                    <SPLIT distance="1100" swimtime="00:12:10.75" />
                    <SPLIT distance="1200" swimtime="00:13:19.96" />
                    <SPLIT distance="1300" swimtime="00:14:29.26" />
                    <SPLIT distance="1400" swimtime="00:15:35.87" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="108" eventid="15" swimtime="00:01:54.22" lane="2" heatid="15009">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:53.63" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="109" eventid="17" swimtime="00:08:26.70" lane="5" heatid="17005">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:57.81" />
                    <SPLIT distance="200" swimtime="00:02:01.10" />
                    <SPLIT distance="300" swimtime="00:03:07.13" />
                    <SPLIT distance="400" swimtime="00:04:11.26" />
                    <SPLIT distance="500" swimtime="00:05:16.41" />
                    <SPLIT distance="600" swimtime="00:06:21.89" />
                    <SPLIT distance="700" swimtime="00:07:26.27" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="110" eventid="31" swimtime="00:00:51.81" lane="6" heatid="31012" />
                <RESULT resultid="111" eventid="33" swimtime="00:04:04.35" lane="3" heatid="33006">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:57.75" />
                    <SPLIT distance="200" swimtime="00:02:00.93" />
                    <SPLIT distance="300" swimtime="00:03:03.80" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="41" birthdate="2009-01-01" gender="M" lastname="Blaszczyk" firstname="Leonard" license="0">
              <RESULTS>
                <RESULT resultid="112" eventid="2" swimtime="00:00:25.81" lane="8" heatid="2003" />
                <RESULT resultid="113" eventid="16" swimtime="00:02:09.37" lane="8" heatid="16003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:01.91" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="114" eventid="32" swimtime="00:00:57.50" lane="2" heatid="32003" />
                <RESULT resultid="115" eventid="34" swimtime="00:04:42.06" lane="1" heatid="34003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:06.03" />
                    <SPLIT distance="200" swimtime="00:02:19.10" />
                    <SPLIT distance="300" swimtime="00:03:33.38" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="42" birthdate="1997-01-01" gender="F" lastname="Walter" firstname="Lisa" license="0">
              <RESULTS>
                <RESULT resultid="116" eventid="3" swimtime="00:16:28.86" lane="8" heatid="3002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:58.70" />
                    <SPLIT distance="200" swimtime="00:02:02.74" />
                    <SPLIT distance="300" swimtime="00:03:07.79" />
                    <SPLIT distance="400" swimtime="00:04:14.02" />
                    <SPLIT distance="500" swimtime="00:05:20.69" />
                    <SPLIT distance="600" swimtime="00:06:27.39" />
                    <SPLIT distance="700" swimtime="00:07:33.87" />
                    <SPLIT distance="800" swimtime="00:08:41.03" />
                    <SPLIT distance="900" swimtime="00:09:47.48" />
                    <SPLIT distance="1000" swimtime="00:10:55.19" />
                    <SPLIT distance="1100" swimtime="00:12:03.20" />
                    <SPLIT distance="1200" swimtime="00:13:11.58" />
                    <SPLIT distance="1300" swimtime="00:14:19.25" />
                    <SPLIT distance="1400" swimtime="00:15:24.76" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="117" eventid="15" swimtime="00:01:56.46" lane="6" heatid="15007">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:54.52" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="118" eventid="17" swimtime="00:08:32.86" lane="7" heatid="17004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:59.06" />
                    <SPLIT distance="200" swimtime="00:02:03.22" />
                    <SPLIT distance="300" swimtime="00:03:07.25" />
                    <SPLIT distance="400" swimtime="00:04:13.02" />
                    <SPLIT distance="500" swimtime="00:05:18.32" />
                    <SPLIT distance="600" swimtime="00:06:24.49" />
                    <SPLIT distance="700" swimtime="00:07:29.82" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="119" eventid="31" swimtime="00:00:54.64" lane="2" heatid="31009" />
                <RESULT resultid="120" eventid="33" swimtime="00:04:16.96" lane="5" heatid="33005">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:00.10" />
                    <SPLIT distance="200" swimtime="00:02:06.25" />
                    <SPLIT distance="300" swimtime="00:03:12.34" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="43" birthdate="2008-01-01" gender="M" lastname="Funke" firstname="Paul" license="0">
              <RESULTS>
                <RESULT resultid="121" eventid="2" swimtime="00:00:22.87" lane="2" heatid="2006" />
                <RESULT resultid="122" eventid="10" swimtime="00:16:55.72" lane="8" heatid="10001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:00.52" />
                    <SPLIT distance="200" swimtime="00:02:08.04" />
                    <SPLIT distance="300" swimtime="00:03:16.27" />
                    <SPLIT distance="400" swimtime="00:04:24.72" />
                    <SPLIT distance="500" swimtime="00:05:33.38" />
                    <SPLIT distance="600" swimtime="00:06:42.67" />
                    <SPLIT distance="700" swimtime="00:07:52.49" />
                    <SPLIT distance="800" swimtime="00:09:03.15" />
                    <SPLIT distance="900" swimtime="00:10:13.38" />
                    <SPLIT distance="1000" swimtime="00:11:23.95" />
                    <SPLIT distance="1100" swimtime="00:12:33.74" />
                    <SPLIT distance="1200" swimtime="00:13:40.69" />
                    <SPLIT distance="1300" swimtime="00:14:47.90" />
                    <SPLIT distance="1400" swimtime="00:15:52.88" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="123" eventid="14" swimtime="00:00:55.55" lane="4" heatid="14001" />
                <RESULT resultid="124" eventid="16" swimtime="00:01:56.31" lane="3" heatid="16005">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:56.66" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="125" eventid="18" swimtime="00:08:46.36" lane="3" heatid="18003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:00.51" />
                    <SPLIT distance="200" swimtime="00:02:07.32" />
                    <SPLIT distance="300" swimtime="00:03:15.33" />
                    <SPLIT distance="400" swimtime="00:04:23.30" />
                    <SPLIT distance="500" swimtime="00:05:31.22" />
                    <SPLIT distance="600" swimtime="00:06:38.65" />
                    <SPLIT distance="700" swimtime="00:07:44.37" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="44" birthdate="2009-01-01" gender="M" lastname="Moritz" firstname="Silas" license="0">
              <RESULTS>
                <RESULT resultid="126" eventid="2" swimtime="00:00:25.22" lane="1" heatid="2005" />
                <RESULT resultid="127" eventid="4" swimtime="00:18:58.10" lane="5" heatid="4001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:07.13" />
                    <SPLIT distance="200" swimtime="00:02:21.75" />
                    <SPLIT distance="300" swimtime="00:03:38.68" />
                    <SPLIT distance="400" swimtime="00:04:55.10" />
                    <SPLIT distance="500" swimtime="00:06:11.51" />
                    <SPLIT distance="600" swimtime="00:07:27.84" />
                    <SPLIT distance="700" swimtime="00:08:45.10" />
                    <SPLIT distance="800" swimtime="00:10:01.55" />
                    <SPLIT distance="900" swimtime="00:11:15.86" />
                    <SPLIT distance="1000" swimtime="00:12:32.09" />
                    <SPLIT distance="1100" swimtime="00:13:49.95" />
                    <SPLIT distance="1200" swimtime="00:15:09.80" />
                    <SPLIT distance="1300" swimtime="00:16:27.60" />
                    <SPLIT distance="1400" swimtime="00:17:44.77" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="128" eventid="16" swimtime="00:02:08.51" lane="2" heatid="16004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:02.15" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="129" eventid="18" swimtime="00:09:32.10" lane="6" heatid="18002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:07.95" />
                    <SPLIT distance="200" swimtime="00:02:21.91" />
                    <SPLIT distance="300" swimtime="00:03:37.30" />
                    <SPLIT distance="400" swimtime="00:04:50.24" />
                    <SPLIT distance="500" swimtime="00:06:02.63" />
                    <SPLIT distance="600" swimtime="00:07:16.26" />
                    <SPLIT distance="700" swimtime="00:08:27.98" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="130" eventid="32" swimtime="00:00:55.71" lane="2" heatid="32005" />
                <RESULT resultid="131" eventid="34" swimtime="00:04:30.70" lane="3" heatid="34003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:02.74" />
                    <SPLIT distance="200" swimtime="00:02:14.71" />
                    <SPLIT distance="300" swimtime="00:03:26.46" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="132" eventid="38" swimtime="00:00:23.80" lane="2" heatid="38003" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY number="1" gender="M" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="89" eventid="49" swimtime="00:03:43.54" lane="4" heatid="49001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:50.30" />
                    <SPLIT distance="200" swimtime="00:01:48.91" />
                    <SPLIT distance="300" swimtime="00:02:45.33" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="39" number="1" />
                    <RELAYPOSITION athleteid="44" number="2" />
                    <RELAYPOSITION athleteid="41" number="3" />
                    <RELAYPOSITION athleteid="38" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" gender="M" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="90" eventid="12" swimtime="00:08:31.78" lane="1" heatid="12002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:55.54" />
                    <SPLIT distance="200" swimtime="00:01:57.51" />
                    <SPLIT distance="300" swimtime="00:02:57.80" />
                    <SPLIT distance="400" swimtime="00:04:06.61" />
                    <SPLIT distance="500" swimtime="00:05:07.06" />
                    <SPLIT distance="600" swimtime="00:06:15.67" />
                    <SPLIT distance="700" swimtime="00:07:17.65" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="43" number="1" />
                    <RELAYPOSITION athleteid="41" number="2" />
                    <RELAYPOSITION athleteid="44" number="3" />
                    <RELAYPOSITION athleteid="38" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" gender="X" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="91" eventid="30" swimtime="00:01:33.40" lane="8" heatid="30003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:48.38" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="43" number="1" />
                    <RELAYPOSITION athleteid="42" number="2" />
                    <RELAYPOSITION athleteid="40" number="3" />
                    <RELAYPOSITION athleteid="39" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB name="COCHTANKLUB Zdar nad Sazavou" nation="CZE" region="0" code="0">
          <ATHLETES>
            <ATHLETE athleteid="54" birthdate="2007-01-01" gender="M" lastname="Styl" firstname="Alan" license="1584">
              <RESULTS>
                <RESULT resultid="165" eventid="6" swimtime="00:00:48.26" lane="2" heatid="6004" />
                <RESULT resultid="163" eventid="14" swimtime="00:00:42.29" lane="2" heatid="14004" />
                <RESULT resultid="164" eventid="32" swimtime="00:00:42.24" lane="2" heatid="32010" />
                <RESULT resultid="166" eventid="40" swimtime="00:00:21.54" lane="3" heatid="40004" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="55" birthdate="2009-01-01" gender="M" lastname="Svoboda" firstname="Jakub" license="1791">
              <RESULTS>
                <RESULT resultid="169" eventid="6" swimtime="00:00:48.98" lane="1" heatid="6004" />
                <RESULT resultid="167" eventid="14" swimtime="00:00:42.65" lane="8" heatid="14005" />
                <RESULT resultid="168" eventid="32" swimtime="00:00:42.31" lane="2" heatid="32012" />
                <RESULT resultid="170" eventid="40" swimtime="00:00:22.54" lane="7" heatid="40004" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="56" birthdate="2008-01-01" gender="F" lastname="Kralickova" firstname="Veronika" license="1439">
              <RESULTS>
                <RESULT resultid="171" eventid="1" swimtime="00:00:21.88" lane="4" heatid="1012" />
                <RESULT resultid="172" eventid="25" swimtime="00:07:32.74" lane="6" heatid="25001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:51.38" />
                    <SPLIT distance="200" swimtime="00:01:47.12" />
                    <SPLIT distance="300" swimtime="00:02:43.82" />
                    <SPLIT distance="400" swimtime="00:03:41.39" />
                    <SPLIT distance="500" swimtime="00:04:39.46" />
                    <SPLIT distance="600" swimtime="00:05:37.93" />
                    <SPLIT distance="700" swimtime="00:06:36.38" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="173" eventid="43" swimtime="00:03:38.78" lane="1" heatid="43001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:49.88" />
                    <SPLIT distance="200" swimtime="00:01:46.09" />
                    <SPLIT distance="300" swimtime="00:02:43.62" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="DJK - VfR Mülheim Saarn" nation="GER" region="28" code="8006000">
          <ATHLETES>
            <ATHLETE athleteid="3" birthdate="1990-01-01" gender="F" lastname="Steenken" firstname="Caroline" license="0">
              <RESULTS>
                <RESULT resultid="3" eventid="1" swimtime="00:00:22.89" lane="3" heatid="1008" />
                <RESULT resultid="4" eventid="13" swimtime="00:00:48.32" lane="1" heatid="13004" />
                <RESULT resultid="5" eventid="15" swimtime="00:01:50.75" lane="1" heatid="15008">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:53.07" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="6" eventid="17" swimtime="00:08:22.65" lane="3" heatid="17003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:58.26" />
                    <SPLIT distance="200" swimtime="00:02:02.06" />
                    <SPLIT distance="300" swimtime="00:03:07.13" />
                    <SPLIT distance="400" swimtime="00:04:12.16" />
                    <SPLIT distance="500" swimtime="00:05:16.41" />
                    <SPLIT distance="600" swimtime="00:06:20.54" />
                    <SPLIT distance="700" swimtime="00:07:23.74" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="7" eventid="31" swimtime="00:00:50.47" lane="5" heatid="31010" />
                <RESULT resultid="8" eventid="33" swimtime="00:04:01.57" lane="4" heatid="33004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:57.43" />
                    <SPLIT distance="200" swimtime="00:01:59.52" />
                    <SPLIT distance="300" swimtime="00:03:02.61" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="4" birthdate="1963-01-01" gender="M" lastname="Venohr" firstname="Heiko" license="0">
              <RESULTS>
                <RESULT resultid="9" eventid="2" swimtime="00:00:21.82" lane="7" heatid="2007" />
                <RESULT resultid="17" eventid="6" swimtime="00:00:55.17" lane="8" heatid="6003" />
                <RESULT resultid="10" eventid="14" swimtime="00:00:43.14" lane="7" heatid="14006" />
                <RESULT resultid="11" eventid="16" swimtime="00:01:49.56" lane="6" heatid="16005">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:53.40" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="12" eventid="18" swimtime="00:08:28.78" lane="5" heatid="18002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:00.08" />
                    <SPLIT distance="200" swimtime="00:02:04.87" />
                    <SPLIT distance="300" swimtime="00:03:10.14" />
                    <SPLIT distance="400" swimtime="00:04:15.21" />
                    <SPLIT distance="500" swimtime="00:05:20.82" />
                    <SPLIT distance="600" swimtime="00:06:25.04" />
                    <SPLIT distance="700" swimtime="00:07:29.27" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="13" eventid="20" swimtime="00:03:47.56" lane="3" heatid="20002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:54.59" />
                    <SPLIT distance="200" swimtime="00:01:51.66" />
                    <SPLIT distance="300" swimtime="00:02:51.38" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="14" eventid="32" swimtime="00:00:51.08" lane="3" heatid="32007" />
                <RESULT resultid="15" eventid="34" swimtime="00:03:55.45" lane="3" heatid="34005">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:56.60" />
                    <SPLIT distance="200" swimtime="00:01:57.53" />
                    <SPLIT distance="300" swimtime="00:02:58.48" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="16" eventid="38" swimtime="00:00:18.49" lane="4" heatid="38006" />
                <RESULT resultid="18" eventid="40" swimtime="00:00:25.68" lane="6" heatid="40002" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="5" birthdate="2005-01-01" gender="M" lastname="Bieler" firstname="Phil Jason" license="0">
              <RESULTS>
                <RESULT resultid="19" eventid="2" swimtime="00:00:19.61" lane="8" heatid="2010" />
                <RESULT resultid="20" eventid="10" swimtime="00:13:50.39" lane="5" heatid="10001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:47.61" />
                    <SPLIT distance="200" swimtime="00:01:41.53" />
                    <SPLIT distance="300" swimtime="00:02:36.29" />
                    <SPLIT distance="400" swimtime="00:03:32.06" />
                    <SPLIT distance="500" swimtime="00:04:27.75" />
                    <SPLIT distance="600" swimtime="00:05:24.59" />
                    <SPLIT distance="700" swimtime="00:06:20.93" />
                    <SPLIT distance="800" swimtime="00:07:17.86" />
                    <SPLIT distance="900" swimtime="00:08:15.26" />
                    <SPLIT distance="1000" swimtime="00:09:12.29" />
                    <SPLIT distance="1100" swimtime="00:10:08.67" />
                    <SPLIT distance="1200" swimtime="00:11:06.32" />
                    <SPLIT distance="1300" swimtime="00:12:01.75" />
                    <SPLIT distance="1400" swimtime="00:12:56.62" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="21" eventid="14" swimtime="00:00:39.58" lane="3" heatid="14004" />
                <RESULT resultid="1501" eventid="22" status="WDR" swimtime="00:00:00.00" lane="0" heatid="22000" />
                <RESULT resultid="22" eventid="26" swimtime="00:07:09.11" lane="5" heatid="26001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:46.47" />
                    <SPLIT distance="200" swimtime="00:01:40.63" />
                    <SPLIT distance="300" swimtime="00:02:35.14" />
                    <SPLIT distance="400" swimtime="00:03:30.14" />
                    <SPLIT distance="500" swimtime="00:04:25.45" />
                    <SPLIT distance="600" swimtime="00:05:20.52" />
                    <SPLIT distance="700" swimtime="00:06:15.97" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="23" eventid="28" swimtime="00:03:13.08" lane="5" heatid="28001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:44.19" />
                    <SPLIT distance="200" swimtime="00:01:34.42" />
                    <SPLIT distance="300" swimtime="00:02:26.22" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="24" eventid="32" swimtime="00:00:42.13" lane="2" heatid="32011" />
                <RESULT resultid="25" eventid="44" swimtime="00:03:24.34" lane="3" heatid="44001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:46.32" />
                    <SPLIT distance="200" swimtime="00:01:39.39" />
                    <SPLIT distance="300" swimtime="00:02:33.69" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="6" birthdate="1977-01-01" gender="F" lastname="Häßler" firstname="Sandra" license="0">
              <RESULTS>
                <RESULT resultid="26" eventid="1" swimtime="00:00:25.11" lane="7" heatid="1006" />
                <RESULT resultid="27" eventid="13" swimtime="00:00:46.66" lane="7" heatid="13007" />
                <RESULT resultid="28" eventid="17" swimtime="00:08:45.95" lane="5" heatid="17003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:00.38" />
                    <SPLIT distance="200" swimtime="00:02:05.17" />
                    <SPLIT distance="300" swimtime="00:03:11.12" />
                    <SPLIT distance="400" swimtime="00:04:17.42" />
                    <SPLIT distance="500" swimtime="00:05:24.05" />
                    <SPLIT distance="600" swimtime="00:06:32.12" />
                    <SPLIT distance="700" swimtime="00:07:40.19" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="29" eventid="19" swimtime="00:03:45.55" lane="1" heatid="19002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:52.71" />
                    <SPLIT distance="200" swimtime="00:01:49.43" />
                    <SPLIT distance="300" swimtime="00:02:48.40" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="30" eventid="33" swimtime="00:04:13.19" lane="4" heatid="33005">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:59.11" />
                    <SPLIT distance="200" swimtime="00:02:02.84" />
                    <SPLIT distance="300" swimtime="00:03:08.79" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="31" eventid="37" swimtime="00:00:21.30" lane="2" heatid="37004" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="7" birthdate="1984-01-01" gender="M" lastname="Link" firstname="Sebastian" license="0">
              <RESULTS>
                <RESULT resultid="32" eventid="2" swimtime="00:00:24.12" lane="4" heatid="2006" />
                <RESULT resultid="37" eventid="6" swimtime="00:00:53.94" lane="8" heatid="6004" />
                <RESULT resultid="33" eventid="16" swimtime="00:01:57.42" lane="1" heatid="16005">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:57.27" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="34" eventid="18" swimtime="00:09:07.18" lane="3" heatid="18002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:01.43" />
                    <SPLIT distance="200" swimtime="00:02:10.96" />
                    <SPLIT distance="300" swimtime="00:03:22.53" />
                    <SPLIT distance="400" swimtime="00:04:34.12" />
                    <SPLIT distance="500" swimtime="00:05:44.67" />
                    <SPLIT distance="600" swimtime="00:06:54.99" />
                    <SPLIT distance="700" swimtime="00:08:04.06" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="35" eventid="32" swimtime="00:00:52.24" lane="1" heatid="32006" />
                <RESULT resultid="36" eventid="34" swimtime="00:04:15.16" lane="2" heatid="34004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:00.07" />
                    <SPLIT distance="200" swimtime="00:02:07.55" />
                    <SPLIT distance="300" swimtime="00:03:15.40" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="38" eventid="40" swimtime="00:00:24.91" lane="2" heatid="40004" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="8" birthdate="2010-01-01" gender="F" lastname="Lazarenko" firstname="Valeria" license="0">
              <RESULTS>
                <RESULT resultid="39" eventid="1" swimtime="00:00:23.16" lane="2" heatid="1010" />
                <RESULT resultid="40" eventid="13" swimtime="00:00:47.15" lane="1" heatid="13006" />
                <RESULT resultid="41" eventid="17" swimtime="00:08:24.00" lane="1" heatid="17004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:56.54" />
                    <SPLIT distance="200" swimtime="00:01:59.78" />
                    <SPLIT distance="300" swimtime="00:03:03.68" />
                    <SPLIT distance="400" swimtime="00:04:08.66" />
                    <SPLIT distance="500" swimtime="00:05:14.17" />
                    <SPLIT distance="600" swimtime="00:06:19.87" />
                    <SPLIT distance="700" swimtime="00:07:23.91" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="42" eventid="19" status="DSQ" swimtime="00:04:06.20" lane="5" heatid="19001" comment="Falscher Start.">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:53.75" />
                    <SPLIT distance="200" swimtime="00:01:57.95" />
                    <SPLIT distance="300" swimtime="00:03:03.48" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="43" eventid="31" swimtime="00:00:51.66" lane="7" heatid="31012" />
                <RESULT resultid="44" eventid="33" swimtime="00:04:05.64" lane="2" heatid="33006">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:58.26" />
                    <SPLIT distance="200" swimtime="00:02:02.15" />
                    <SPLIT distance="300" swimtime="00:03:05.69" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="45" eventid="35" swimtime="00:00:20.81" lane="4" heatid="35002" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY number="15" gender="X" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="1" eventid="29" swimtime="00:01:35.92" lane="4" heatid="29001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:49.58" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="7" number="1" />
                    <RELAYPOSITION athleteid="6" number="2" />
                    <RELAYPOSITION athleteid="4" number="3" />
                    <RELAYPOSITION athleteid="3" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="25" gender="X" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="2" eventid="47" swimtime="00:03:28.76" lane="4" heatid="47001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:52.35" />
                    <SPLIT distance="200" swimtime="00:01:42.61" />
                    <SPLIT distance="300" swimtime="00:02:32.66" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="7" number="1" />
                    <RELAYPOSITION athleteid="3" number="2" />
                    <RELAYPOSITION athleteid="4" number="3" />
                    <RELAYPOSITION athleteid="6" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB name="HSTSG Hamburg" nation="GER" region="23" code="0">
          <ATHLETES>
            <ATHLETE athleteid="196" birthdate="1962-11-22" gender="M" lastname="Bandilla" firstname="Dalk-Ascan" license="0">
              <RESULTS>
                <RESULT resultid="735" eventid="2" swimtime="00:00:26.59" lane="6" heatid="2002" />
                <RESULT resultid="736" eventid="6" swimtime="00:01:00.70" lane="2" heatid="6002" />
                <RESULT resultid="737" eventid="16" swimtime="00:02:18.90" lane="8" heatid="16002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:05.14" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="738" eventid="18" swimtime="00:10:59.24" lane="2" heatid="18001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:12.42" />
                    <SPLIT distance="200" swimtime="00:02:35.64" />
                    <SPLIT distance="300" swimtime="00:03:59.65" />
                    <SPLIT distance="400" swimtime="00:05:25.26" />
                    <SPLIT distance="500" swimtime="00:06:51.66" />
                    <SPLIT distance="600" swimtime="00:08:17.46" />
                    <SPLIT distance="700" swimtime="00:09:42.71" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="739" eventid="32" swimtime="00:00:58.85" lane="4" heatid="32002" />
                <RESULT resultid="740" eventid="34" swimtime="00:05:18.16" lane="3" heatid="34002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:13.20" />
                    <SPLIT distance="200" swimtime="00:02:35.33" />
                    <SPLIT distance="300" swimtime="00:04:00.83" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="741" eventid="40" swimtime="00:00:26.73" lane="3" heatid="40001" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="SC DHfK Leipzig Flossenschwimmen" nation="GER" region="20" code="0">
          <ATHLETES>
            <ATHLETE athleteid="240" birthdate="2001-01-01" gender="F" lastname="Hecke" firstname="Aimee Joy" license="0">
              <RESULTS>
                <RESULT resultid="913" eventid="31" status="DNS" swimtime="00:00:00.00" lane="8" heatid="31016" />
                <RESULT resultid="914" eventid="39" status="DNS" swimtime="00:00:00.00" lane="2" heatid="39004" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="241" birthdate="2008-01-01" gender="M" lastname="Berger" firstname="Alex Michael" license="0">
              <RESULTS>
                <RESULT resultid="915" eventid="2" swimtime="00:00:20.30" lane="7" heatid="2008" />
                <RESULT resultid="916" eventid="16" swimtime="00:01:42.95" lane="1" heatid="16008">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:48.77" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="917" eventid="32" swimtime="00:00:45.81" lane="5" heatid="32008" />
                <RESULT resultid="918" eventid="34" swimtime="00:03:53.10" lane="2" heatid="34006">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:54.75" />
                    <SPLIT distance="200" swimtime="00:01:55.81" />
                    <SPLIT distance="300" swimtime="00:02:57.58" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="919" eventid="38" swimtime="00:00:19.45" lane="1" heatid="38005" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="242" birthdate="2001-01-01" gender="F" lastname="Franke" firstname="Aleyna" license="0">
              <RESULTS>
                <RESULT resultid="920" eventid="31" swimtime="00:00:47.51" lane="7" heatid="31013" />
                <RESULT resultid="921" eventid="37" swimtime="00:00:19.64" lane="2" heatid="37006" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="243" birthdate="2007-01-01" gender="M" lastname="Schoodt" firstname="Ben Joseph" license="2944">
              <RESULTS>
                <RESULT resultid="922" eventid="2" swimtime="00:00:17.77" lane="3" heatid="2011" />
                <RESULT resultid="1417" eventid="8" swimtime="00:00:18.03" lane="7" heatid="8001" />
                <RESULT resultid="923" eventid="16" swimtime="00:01:33.21" lane="3" heatid="16006">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:43.66" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1531" eventid="24" swimtime="00:01:33.52" lane="2" heatid="24001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:44.32" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="924" eventid="32" swimtime="00:00:41.39" lane="6" heatid="32012" />
                <RESULT resultid="926" eventid="38" swimtime="00:00:17.03" lane="3" heatid="38009" />
                <RESULT resultid="925" eventid="44" swimtime="00:03:47.55" lane="1" heatid="44001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:51.21" />
                    <SPLIT distance="200" swimtime="00:01:49.32" />
                    <SPLIT distance="300" swimtime="00:02:49.19" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="244" birthdate="1998-01-01" gender="F" lastname="Gerungan" firstname="Daveena" license="0">
              <RESULTS>
                <RESULT resultid="927" eventid="1" swimtime="00:00:22.27" lane="8" heatid="1014" />
                <RESULT resultid="928" eventid="15" swimtime="00:01:49.31" lane="6" heatid="15009">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:51.10" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="929" eventid="31" swimtime="00:00:46.43" lane="4" heatid="31014" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="245" birthdate="2001-01-01" gender="M" lastname="Gaida" firstname="Duncan" license="0">
              <RESULTS>
                <RESULT resultid="930" eventid="10" swimtime="00:12:54.90" lane="4" heatid="10001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:47.37" />
                    <SPLIT distance="200" swimtime="00:01:37.69" />
                    <SPLIT distance="300" swimtime="00:02:28.59" />
                    <SPLIT distance="400" swimtime="00:03:20.13" />
                    <SPLIT distance="500" swimtime="00:04:12.26" />
                    <SPLIT distance="600" swimtime="00:05:04.53" />
                    <SPLIT distance="700" swimtime="00:05:56.82" />
                    <SPLIT distance="800" swimtime="00:06:49.22" />
                    <SPLIT distance="900" swimtime="00:07:41.72" />
                    <SPLIT distance="1000" swimtime="00:08:34.34" />
                    <SPLIT distance="1100" swimtime="00:09:26.79" />
                    <SPLIT distance="1200" swimtime="00:10:19.75" />
                    <SPLIT distance="1300" swimtime="00:11:12.32" />
                    <SPLIT distance="1400" swimtime="00:12:04.68" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="931" eventid="16" swimtime="00:01:27.78" lane="4" heatid="16006">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:42.94" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1524" eventid="24" status="WDR" swimtime="00:00:00.00" lane="0" heatid="24000" />
                <RESULT resultid="932" eventid="26" swimtime="00:06:39.30" lane="4" heatid="26001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:46.62" />
                    <SPLIT distance="200" swimtime="00:01:36.38" />
                    <SPLIT distance="300" swimtime="00:02:26.64" />
                    <SPLIT distance="400" swimtime="00:03:17.51" />
                    <SPLIT distance="500" swimtime="00:04:08.47" />
                    <SPLIT distance="600" swimtime="00:04:59.70" />
                    <SPLIT distance="700" swimtime="00:05:50.48" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="933" eventid="44" swimtime="00:03:11.88" lane="4" heatid="44001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:45.36" />
                    <SPLIT distance="200" swimtime="00:01:34.32" />
                    <SPLIT distance="300" swimtime="00:02:23.56" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="246" birthdate="2007-01-01" gender="F" lastname="Hempler" firstname="Emily" license="0">
              <RESULTS>
                <RESULT resultid="934" eventid="9" swimtime="00:14:25.03" lane="5" heatid="9001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:52.48" />
                    <SPLIT distance="200" swimtime="00:01:48.16" />
                    <SPLIT distance="300" swimtime="00:02:45.12" />
                    <SPLIT distance="400" swimtime="00:03:43.13" />
                    <SPLIT distance="500" swimtime="00:04:41.18" />
                    <SPLIT distance="600" swimtime="00:05:39.51" />
                    <SPLIT distance="700" swimtime="00:06:38.09" />
                    <SPLIT distance="800" swimtime="00:07:36.89" />
                    <SPLIT distance="900" swimtime="00:08:35.43" />
                    <SPLIT distance="1000" swimtime="00:09:34.11" />
                    <SPLIT distance="1100" swimtime="00:10:32.58" />
                    <SPLIT distance="1200" swimtime="00:11:31.41" />
                    <SPLIT distance="1300" swimtime="00:12:29.81" />
                    <SPLIT distance="1400" swimtime="00:13:27.94" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="935" eventid="15" swimtime="00:01:41.19" lane="2" heatid="15012">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:48.32" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1513" eventid="23" status="WDR" swimtime="00:00:00.00" lane="0" heatid="23000" />
                <RESULT resultid="936" eventid="25" swimtime="00:07:30.13" lane="5" heatid="25001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:50.99" />
                    <SPLIT distance="200" swimtime="00:01:46.71" />
                    <SPLIT distance="300" swimtime="00:02:43.76" />
                    <SPLIT distance="400" swimtime="00:03:41.52" />
                    <SPLIT distance="500" swimtime="00:04:39.92" />
                    <SPLIT distance="600" swimtime="00:05:38.01" />
                    <SPLIT distance="700" swimtime="00:06:34.67" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="937" eventid="31" swimtime="00:00:45.05" lane="4" heatid="31013" />
                <RESULT resultid="938" eventid="43" swimtime="00:03:35.44" lane="3" heatid="43001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:49.36" />
                    <SPLIT distance="200" swimtime="00:01:43.90" />
                    <SPLIT distance="300" swimtime="00:02:40.23" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="247" birthdate="1999-01-01" gender="M" lastname="Wahlstadt" firstname="Felix" license="267">
              <RESULTS>
                <RESULT resultid="939" eventid="2" swimtime="00:00:17.89" lane="5" heatid="2011" />
                <RESULT resultid="1418" eventid="8" swimtime="00:00:17.74" lane="1" heatid="8001" />
                <RESULT resultid="940" eventid="16" swimtime="00:01:31.27" lane="3" heatid="16008">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:43.51" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1530" eventid="24" swimtime="00:01:29.72" lane="6" heatid="24001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:43.04" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="941" eventid="32" swimtime="00:00:41.56" lane="3" heatid="32011" />
                <RESULT resultid="942" eventid="44" swimtime="00:03:21.86" lane="2" heatid="44001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:45.76" />
                    <SPLIT distance="200" swimtime="00:01:35.84" />
                    <SPLIT distance="300" swimtime="00:02:28.13" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="248" birthdate="2011-01-01" gender="F" lastname="Hau" firstname="Hannah" license="0">
              <RESULTS>
                <RESULT resultid="943" eventid="1" swimtime="00:00:28.84" lane="5" heatid="1001" />
                <RESULT resultid="944" eventid="15" swimtime="00:02:20.94" lane="4" heatid="15001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:04.81" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="945" eventid="31" swimtime="00:01:02.06" lane="2" heatid="31002" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="249" birthdate="2001-01-01" gender="M" lastname="Mörstedt" firstname="Justus" license="0">
              <RESULTS>
                <RESULT resultid="946" eventid="14" swimtime="00:00:33.87" lane="4" heatid="14005" />
                <RESULT resultid="947" eventid="16" swimtime="00:01:27.05" lane="4" heatid="16008">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:41.54" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1504" eventid="22" swimtime="00:00:32.37" lane="4" heatid="22001" />
                <RESULT resultid="1527" eventid="24" swimtime="00:01:21.26" lane="4" heatid="24001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:39.11" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="948" eventid="32" swimtime="00:00:36.89" lane="4" heatid="32011" />
                <RESULT resultid="949" eventid="38" swimtime="00:00:14.94" lane="4" heatid="38008" />
                <RESULT resultid="1543" eventid="42" swimtime="00:00:34.73" lane="4" heatid="42001" />
                <RESULT resultid="1561" eventid="46" swimtime="00:00:14.49" lane="3" heatid="46001" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="250" birthdate="1997-01-01" gender="F" lastname="Vos" firstname="Katharina" license="0">
              <RESULTS>
                <RESULT resultid="950" eventid="1" swimtime="00:00:20.92" lane="6" heatid="1015" />
                <RESULT resultid="951" eventid="39" swimtime="00:00:24.01" lane="5" heatid="39004" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="251" birthdate="2008-01-01" gender="F" lastname="Säbisch" firstname="Kyra" license="0">
              <RESULTS>
                <RESULT resultid="952" eventid="1" swimtime="00:00:21.10" lane="8" heatid="1013" />
                <RESULT resultid="953" eventid="15" swimtime="00:01:49.11" lane="3" heatid="15007">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:52.21" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="954" eventid="31" swimtime="00:00:47.47" lane="6" heatid="31010" />
                <RESULT resultid="955" eventid="37" swimtime="00:00:19.36" lane="1" heatid="37005" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="252" birthdate="2007-01-01" gender="F" lastname="Holtz" firstname="Leonie-Florentine" license="2947">
              <RESULTS>
                <RESULT resultid="956" eventid="1" swimtime="00:00:24.04" lane="8" heatid="1010" />
                <RESULT resultid="957" eventid="13" swimtime="00:00:51.53" lane="4" heatid="13004" />
                <RESULT resultid="958" eventid="31" swimtime="00:00:55.31" lane="5" heatid="31009" />
                <RESULT resultid="959" eventid="37" swimtime="00:00:22.68" lane="4" heatid="37002" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="253" birthdate="2008-01-01" gender="F" lastname="Horenok" firstname="Maiia" license="0">
              <RESULTS>
                <RESULT resultid="960" eventid="1" swimtime="00:00:19.66" lane="5" heatid="1015" />
                <RESULT resultid="1408" eventid="7" swimtime="00:00:18.97" lane="2" heatid="7001" />
                <RESULT resultid="961" eventid="13" swimtime="00:00:41.53" lane="5" heatid="13005" />
                <RESULT resultid="962" eventid="15" swimtime="00:01:39.11" lane="5" heatid="15010">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:47.89" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1498" eventid="21" swimtime="00:00:42.07" lane="7" heatid="21001" />
                <RESULT resultid="1519" eventid="23" swimtime="00:01:39.24" lane="7" heatid="23001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:47.43" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="963" eventid="31" swimtime="00:00:43.91" lane="5" heatid="31017" />
                <RESULT resultid="964" eventid="37" swimtime="00:00:17.68" lane="4" heatid="37007" />
                <RESULT resultid="1541" eventid="41" swimtime="00:00:42.85" lane="1" heatid="41001" />
                <RESULT resultid="1552" eventid="45" swimtime="00:00:17.59" lane="5" heatid="45001" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="254" birthdate="1994-01-01" gender="M" lastname="Poschart" firstname="Max" license="0">
              <RESULTS>
                <RESULT resultid="965" eventid="2" swimtime="00:00:16.16" lane="4" heatid="2011" />
                <RESULT resultid="1413" eventid="8" swimtime="00:00:15.28" lane="5" heatid="8001" />
                <RESULT resultid="966" eventid="14" swimtime="00:00:37.67" lane="4" heatid="14006" />
                <RESULT resultid="967" eventid="16" swimtime="00:01:20.94" lane="4" heatid="16007">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:39.26" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1507" eventid="22" swimtime="00:00:32.39" lane="6" heatid="22001" />
                <RESULT resultid="1525" eventid="24" status="WDR" swimtime="00:00:00.00" lane="0" heatid="24000" />
                <RESULT resultid="968" eventid="32" swimtime="00:00:39.07" lane="4" heatid="32012" />
                <RESULT resultid="969" eventid="38" swimtime="00:00:14.23" lane="4" heatid="38009" />
                <RESULT resultid="1545" eventid="42" swimtime="00:00:34.08" lane="3" heatid="42001" />
                <RESULT resultid="1559" eventid="46" swimtime="00:00:14.41" lane="4" heatid="46001" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="255" birthdate="2009-01-01" gender="M" lastname="Batiuk" firstname="Mykyta" license="0">
              <RESULTS>
                <RESULT resultid="970" eventid="2" swimtime="00:00:19.25" lane="7" heatid="2009" />
                <RESULT resultid="971" eventid="32" swimtime="00:00:46.12" lane="1" heatid="32009" />
                <RESULT resultid="972" eventid="38" swimtime="00:00:17.81" lane="6" heatid="38006" />
                <RESULT resultid="973" eventid="40" swimtime="00:00:23.66" lane="2" heatid="40003" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="256" birthdate="2004-01-01" gender="F" lastname="Barthel" firstname="Nadja" license="0">
              <RESULTS>
                <RESULT resultid="974" eventid="1" swimtime="00:00:19.13" lane="4" heatid="1014" />
                <RESULT resultid="1405" eventid="7" swimtime="00:00:19.47" lane="5" heatid="7001" />
                <RESULT resultid="975" eventid="15" swimtime="00:01:36.52" lane="4" heatid="15010">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:46.26" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1517" eventid="23" swimtime="00:01:35.51" lane="6" heatid="23001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:46.02" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="976" eventid="31" swimtime="00:00:42.51" lane="4" heatid="31016" />
                <RESULT resultid="977" eventid="39" status="DNS" swimtime="00:00:00.00" lane="6" heatid="39004" />
                <RESULT resultid="1535" eventid="41" swimtime="00:00:42.58" lane="4" heatid="41001" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="257" birthdate="2010-01-01" gender="F" lastname="Horenok" firstname="Polina" license="0">
              <RESULTS>
                <RESULT resultid="978" eventid="1" swimtime="00:00:25.00" lane="2" heatid="1005" />
                <RESULT resultid="979" eventid="13" swimtime="00:01:00.50" lane="6" heatid="13001" />
                <RESULT resultid="980" eventid="31" swimtime="00:00:57.88" lane="8" heatid="31006" />
                <RESULT resultid="981" eventid="35" swimtime="00:00:25.95" lane="8" heatid="35002" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="258" birthdate="2008-01-01" gender="F" lastname="Kulchytska" firstname="Polina" license="0">
              <RESULTS>
                <RESULT resultid="982" eventid="9" swimtime="00:15:37.70" lane="6" heatid="9001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:56.36" />
                    <SPLIT distance="200" swimtime="00:01:59.48" />
                    <SPLIT distance="300" swimtime="00:03:02.49" />
                    <SPLIT distance="400" swimtime="00:04:05.85" />
                    <SPLIT distance="500" swimtime="00:05:09.81" />
                    <SPLIT distance="600" swimtime="00:06:14.39" />
                    <SPLIT distance="700" swimtime="00:07:16.45" />
                    <SPLIT distance="800" swimtime="00:08:20.97" />
                    <SPLIT distance="900" swimtime="00:09:23.96" />
                    <SPLIT distance="1000" swimtime="00:10:28.32" />
                    <SPLIT distance="1100" swimtime="00:11:33.19" />
                    <SPLIT distance="1200" swimtime="00:12:37.01" />
                    <SPLIT distance="1300" swimtime="00:13:38.68" />
                    <SPLIT distance="1400" swimtime="00:14:39.16" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="983" eventid="13" swimtime="00:00:44.59" lane="3" heatid="13006" />
                <RESULT resultid="984" eventid="17" swimtime="00:08:08.73" lane="4" heatid="17005">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:58.79" />
                    <SPLIT distance="200" swimtime="00:02:01.16" />
                    <SPLIT distance="300" swimtime="00:03:03.91" />
                    <SPLIT distance="400" swimtime="00:04:05.71" />
                    <SPLIT distance="500" swimtime="00:05:08.86" />
                    <SPLIT distance="600" swimtime="00:06:10.27" />
                    <SPLIT distance="700" swimtime="00:07:10.81" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="985" eventid="31" swimtime="00:00:48.83" lane="6" heatid="31013" />
                <RESULT resultid="986" eventid="33" swimtime="00:03:55.75" lane="4" heatid="33006">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:55.89" />
                    <SPLIT distance="200" swimtime="00:01:57.35" />
                    <SPLIT distance="300" swimtime="00:02:58.11" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="259" birthdate="1996-01-01" gender="M" lastname="Zeuner" firstname="Sidney" license="0">
              <RESULTS>
                <RESULT resultid="987" eventid="2" swimtime="00:00:17.16" lane="5" heatid="2009" />
                <RESULT resultid="1415" eventid="8" swimtime="00:00:16.74" lane="6" heatid="8001" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="260" birthdate="1998-01-01" gender="F" lastname="Niemann" firstname="Sophie" license="0">
              <RESULTS>
                <RESULT resultid="988" eventid="31" swimtime="00:00:45.27" lane="7" heatid="31015" />
                <RESULT resultid="989" eventid="37" swimtime="00:00:18.72" lane="6" heatid="37006" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="262" birthdate="1958-01-01" gender="F" lastname="Hirschfeldt" firstname="Birgit" license="0">
              <RESULTS>
                <RESULT resultid="992" eventid="1" swimtime="00:00:31.19" lane="1" heatid="1001" />
                <RESULT resultid="994" eventid="5" swimtime="00:01:16.22" lane="5" heatid="5001" />
                <RESULT resultid="993" eventid="31" swimtime="00:01:13.82" lane="3" heatid="31001" />
                <RESULT resultid="995" eventid="39" swimtime="00:00:33.28" lane="2" heatid="39001" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="263" birthdate="1987-01-01" gender="F" lastname="Eckstein" firstname="Diana" license="0">
              <RESULTS>
                <RESULT resultid="996" eventid="1" swimtime="00:00:24.68" lane="7" heatid="1008" />
                <RESULT resultid="998" eventid="5" swimtime="00:01:03.05" lane="2" heatid="5003" />
                <RESULT resultid="997" eventid="31" swimtime="00:00:55.14" lane="1" heatid="31008" />
                <RESULT resultid="999" eventid="39" swimtime="00:00:27.73" lane="7" heatid="39003" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="264" birthdate="1984-01-01" gender="F" lastname="Sapsai" firstname="Iryna" license="0">
              <RESULTS>
                <RESULT resultid="1000" eventid="1" status="DSQ" swimtime="00:00:24.31" lane="6" heatid="1007" comment="Falsche Ausrüstung." />
                <RESULT resultid="1001" eventid="39" swimtime="00:00:27.90" lane="8" heatid="39003" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="265" birthdate="1966-01-01" gender="M" lastname="Weigang" firstname="Mike" license="0">
              <RESULTS>
                <RESULT resultid="1002" eventid="6" swimtime="00:00:57.81" lane="5" heatid="6001" />
                <RESULT resultid="1003" eventid="40" swimtime="00:00:26.28" lane="8" heatid="40002" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="266" birthdate="1978-01-01" gender="M" lastname="Bordag" firstname="Stefan" license="0">
              <RESULTS>
                <RESULT resultid="1375" eventid="2" swimtime="00:00:24.87" lane="2" heatid="2005" />
                <RESULT resultid="1006" eventid="6" swimtime="00:00:58.56" lane="1" heatid="6002" />
                <RESULT resultid="1004" eventid="32" swimtime="00:00:54.23" lane="5" heatid="32004" />
                <RESULT resultid="1005" eventid="38" swimtime="00:00:22.06" lane="3" heatid="38003" />
                <RESULT resultid="1007" eventid="40" swimtime="00:00:26.61" lane="1" heatid="40002" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="267" birthdate="1977-01-01" gender="M" lastname="Nehrdich" firstname="Thomas" license="0">
              <RESULTS>
                <RESULT resultid="1008" eventid="2" swimtime="00:00:20.03" lane="5" heatid="2008" />
                <RESULT resultid="1012" eventid="6" swimtime="00:00:53.20" lane="4" heatid="6003" />
                <RESULT resultid="1009" eventid="16" swimtime="00:01:45.27" lane="8" heatid="16007">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:50.29" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1010" eventid="32" status="DSQ" swimtime="00:00:45.76" lane="3" heatid="32008" comment="Falscher Start." />
                <RESULT resultid="1011" eventid="34" swimtime="00:03:51.05" lane="6" heatid="34006">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:53.03" />
                    <SPLIT distance="200" swimtime="00:01:52.87" />
                    <SPLIT distance="300" swimtime="00:02:54.02" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1013" eventid="40" swimtime="00:00:23.36" lane="6" heatid="40003" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="268" birthdate="1973-01-01" gender="M" lastname="Stelzig" firstname="Torsten" license="0">
              <RESULTS>
                <RESULT resultid="1014" eventid="2" swimtime="00:00:24.50" lane="5" heatid="2004" />
                <RESULT resultid="1017" eventid="6" swimtime="00:00:59.45" lane="8" heatid="6002" />
                <RESULT resultid="1015" eventid="32" swimtime="00:00:55.50" lane="3" heatid="32004" />
                <RESULT resultid="1016" eventid="38" swimtime="00:00:22.50" lane="6" heatid="38003" />
                <RESULT resultid="1018" eventid="40" swimtime="00:00:26.79" lane="4" heatid="40001" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="269" birthdate="1969-01-01" gender="F" lastname="Meier-Mahlo" firstname="Ulrike" license="0">
              <RESULTS>
                <RESULT resultid="1019" eventid="1" swimtime="00:00:24.44" lane="1" heatid="1008" />
                <RESULT resultid="1022" eventid="5" swimtime="00:01:02.01" lane="7" heatid="5003" />
                <RESULT resultid="1020" eventid="31" swimtime="00:00:54.87" lane="3" heatid="31007" />
                <RESULT resultid="1021" eventid="37" swimtime="00:00:22.21" lane="8" heatid="37003" />
                <RESULT resultid="1023" eventid="39" swimtime="00:00:28.20" lane="4" heatid="39002" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="270" birthdate="1967-01-01" gender="M" lastname="Meier" firstname="Wolf-Dieter" license="0">
              <RESULTS>
                <RESULT resultid="1024" eventid="2" swimtime="00:00:22.87" lane="4" heatid="2005" />
                <RESULT resultid="1026" eventid="6" swimtime="00:00:56.63" lane="1" heatid="6003" />
                <RESULT resultid="1025" eventid="34" swimtime="00:04:16.58" lane="3" heatid="34004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:59.45" />
                    <SPLIT distance="200" swimtime="00:02:05.18" />
                    <SPLIT distance="300" swimtime="00:03:12.07" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1027" eventid="40" swimtime="00:00:25.48" lane="8" heatid="40003" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY number="1" gender="M" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="904" eventid="12" swimtime="00:05:40.84" lane="4" heatid="12002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:37.08" />
                    <SPLIT distance="200" swimtime="00:01:21.13" />
                    <SPLIT distance="300" swimtime="00:02:03.08" />
                    <SPLIT distance="400" swimtime="00:02:48.86" />
                    <SPLIT distance="500" swimtime="00:03:31.22" />
                    <SPLIT distance="600" swimtime="00:04:20.42" />
                    <SPLIT distance="700" swimtime="00:04:58.20" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="249" number="1" />
                    <RELAYPOSITION athleteid="245" number="2" />
                    <RELAYPOSITION athleteid="247" number="3" />
                    <RELAYPOSITION athleteid="254" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT resultid="905" eventid="49" swimtime="00:02:29.24" lane="4" heatid="49002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:41.47" />
                    <SPLIT distance="200" swimtime="00:01:15.12" />
                    <SPLIT distance="300" swimtime="00:01:51.21" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="243" number="1" />
                    <RELAYPOSITION athleteid="254" number="2" />
                    <RELAYPOSITION athleteid="249" number="3" />
                    <RELAYPOSITION athleteid="245" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" gender="X" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="906" eventid="30" swimtime="00:01:10.34" lane="4" heatid="30004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:36.67" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="249" number="1" />
                    <RELAYPOSITION athleteid="250" number="2" />
                    <RELAYPOSITION athleteid="254" number="3" />
                    <RELAYPOSITION athleteid="256" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" gender="F" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="907" eventid="11" swimtime="00:06:49.59" lane="3" heatid="11003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:47.25" />
                    <SPLIT distance="200" swimtime="00:01:38.41" />
                    <SPLIT distance="300" swimtime="00:02:25.51" />
                    <SPLIT distance="400" swimtime="00:03:19.80" />
                    <SPLIT distance="500" swimtime="00:04:11.95" />
                    <SPLIT distance="600" swimtime="00:05:12.45" />
                    <SPLIT distance="700" swimtime="00:05:56.35" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="253" number="1" />
                    <RELAYPOSITION athleteid="246" number="2" />
                    <RELAYPOSITION athleteid="251" number="3" />
                    <RELAYPOSITION athleteid="256" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT resultid="908" eventid="48" swimtime="00:02:56.95" lane="3" heatid="48003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:42.85" />
                    <SPLIT distance="200" swimtime="00:01:28.90" />
                    <SPLIT distance="300" swimtime="00:02:12.40" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="256" number="1" />
                    <RELAYPOSITION athleteid="242" number="2" />
                    <RELAYPOSITION athleteid="246" number="3" />
                    <RELAYPOSITION athleteid="260" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="2" gender="F" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="909" eventid="48" swimtime="00:03:19.40" lane="3" heatid="48002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:48.60" />
                    <SPLIT distance="200" swimtime="00:01:32.80" />
                    <SPLIT distance="300" swimtime="00:02:33.49" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="251" number="1" />
                    <RELAYPOSITION athleteid="253" number="2" />
                    <RELAYPOSITION athleteid="248" number="3" />
                    <RELAYPOSITION athleteid="244" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="2" gender="X" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="910" eventid="30" swimtime="00:01:20.62" lane="1" heatid="30004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:38.95" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="243" number="1" />
                    <RELAYPOSITION athleteid="246" number="2" />
                    <RELAYPOSITION athleteid="241" number="3" />
                    <RELAYPOSITION athleteid="251" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="2" gender="F" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="911" eventid="11" swimtime="00:08:19.06" lane="7" heatid="11002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:50.96" />
                    <SPLIT distance="200" swimtime="00:01:49.05" />
                    <SPLIT distance="300" swimtime="00:02:40.77" />
                    <SPLIT distance="400" swimtime="00:03:39.82" />
                    <SPLIT distance="500" swimtime="00:04:41.62" />
                    <SPLIT distance="600" swimtime="00:05:54.26" />
                    <SPLIT distance="700" swimtime="00:07:00.18" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="244" number="1" />
                    <RELAYPOSITION athleteid="258" number="2" />
                    <RELAYPOSITION athleteid="257" number="3" />
                    <RELAYPOSITION athleteid="248" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="3" gender="X" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="912" eventid="30" swimtime="00:01:19.04" lane="7" heatid="30004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:36.10" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="245" number="1" />
                    <RELAYPOSITION athleteid="253" number="2" />
                    <RELAYPOSITION athleteid="247" number="3" />
                    <RELAYPOSITION athleteid="257" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="100" gender="X" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="990" eventid="29" swimtime="00:01:32.65" lane="5" heatid="29001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:49.72" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="263" number="1" />
                    <RELAYPOSITION athleteid="264" number="2" />
                    <RELAYPOSITION athleteid="265" number="3" />
                    <RELAYPOSITION athleteid="267" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT resultid="991" eventid="47" swimtime="00:03:31.07" lane="5" heatid="47001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:56.84" />
                    <SPLIT distance="200" swimtime="00:01:53.30" />
                    <SPLIT distance="300" swimtime="00:02:46.06" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="263" number="1" />
                    <RELAYPOSITION athleteid="269" number="2" />
                    <RELAYPOSITION athleteid="270" number="3" />
                    <RELAYPOSITION athleteid="267" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB name="SC Riesa Sekt Flossenschwimmen" nation="GER" region="20" code="154149">
          <ATHLETES>
            <ATHLETE athleteid="205" birthdate="2011-01-01" gender="F" lastname="Hönisch" firstname="Ida" license="0">
              <RESULTS>
                <RESULT resultid="787" eventid="1" swimtime="00:00:28.98" lane="1" heatid="1002" />
                <RESULT resultid="788" eventid="15" swimtime="00:02:24.17" lane="3" heatid="15002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:08.25" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="789" eventid="31" swimtime="00:01:02.08" lane="3" heatid="31003" />
                <RESULT resultid="790" eventid="33" swimtime="00:05:18.04" lane="8" heatid="33002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:12.38" />
                    <SPLIT distance="200" swimtime="00:02:35.43" />
                    <SPLIT distance="300" swimtime="00:04:00.11" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="206" birthdate="2010-01-01" gender="F" lastname="Berger" firstname="Lene" license="0">
              <RESULTS>
                <RESULT resultid="791" eventid="1" swimtime="00:00:27.07" lane="1" heatid="1004" />
                <RESULT resultid="792" eventid="15" swimtime="00:02:13.06" lane="2" heatid="15004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:01.59" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="793" eventid="31" swimtime="00:00:58.91" lane="1" heatid="31005" />
                <RESULT resultid="794" eventid="33" swimtime="00:04:45.26" lane="4" heatid="33002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:04.75" />
                    <SPLIT distance="200" swimtime="00:02:20.40" />
                    <SPLIT distance="300" swimtime="00:03:34.70" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="207" birthdate="2006-01-01" gender="M" lastname="Loßner" firstname="Niklas" license="0">
              <RESULTS>
                <RESULT resultid="795" eventid="2" swimtime="00:00:15.90" lane="4" heatid="2010" />
                <RESULT resultid="1412" eventid="8" swimtime="00:00:16.09" lane="4" heatid="8001" />
                <RESULT resultid="796" eventid="14" swimtime="00:00:37.58" lane="4" heatid="14004" />
                <RESULT resultid="797" eventid="16" swimtime="00:01:29.77" lane="5" heatid="16007">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:41.16" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1506" eventid="22" swimtime="00:00:33.75" lane="3" heatid="22001" />
                <RESULT resultid="1523" eventid="24" status="WDR" swimtime="00:00:00.00" lane="0" heatid="24000" />
                <RESULT resultid="798" eventid="32" swimtime="00:00:40.48" lane="5" heatid="32012" />
                <RESULT resultid="799" eventid="38" swimtime="00:00:14.36" lane="4" heatid="38007" />
                <RESULT resultid="1549" eventid="42" swimtime="00:00:36.63" lane="1" heatid="42001" />
                <RESULT resultid="1560" eventid="46" swimtime="00:00:14.19" lane="5" heatid="46001" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="SG Dresden (TC)" nation="GER" region="20" code="0">
          <ATHLETES>
            <ATHLETE athleteid="198" birthdate="2005-01-01" gender="F" lastname="Richter" firstname="Franca" license="0">
              <RESULTS>
                <RESULT resultid="744" eventid="1" swimtime="00:00:20.27" lane="6" heatid="1013" />
                <RESULT resultid="745" eventid="13" swimtime="00:00:40.97" lane="4" heatid="13005" />
                <RESULT resultid="746" eventid="15" status="DNS" swimtime="00:00:00.00" lane="3" heatid="15012" />
                <RESULT resultid="1492" eventid="21" status="WDR" swimtime="00:00:00.00" lane="0" heatid="21000" />
                <RESULT resultid="747" eventid="27" status="DNS" swimtime="00:00:00.00" lane="4" heatid="27001" />
                <RESULT resultid="748" eventid="31" status="DNS" swimtime="00:00:00.00" lane="3" heatid="31015" />
                <RESULT resultid="749" eventid="43" status="DNS" swimtime="00:00:00.00" lane="5" heatid="43001" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="199" birthdate="1943-01-01" gender="M" lastname="Pietzsch" firstname="Gerd" license="0">
              <RESULTS>
                <RESULT resultid="750" eventid="2" swimtime="00:00:32.14" lane="5" heatid="2001" />
                <RESULT resultid="752" eventid="16" swimtime="00:02:51.51" lane="5" heatid="16001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:16.84" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="753" eventid="18" swimtime="00:12:38.08" lane="5" heatid="18001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:24.75" />
                    <SPLIT distance="200" swimtime="00:03:03.14" />
                    <SPLIT distance="300" swimtime="00:04:40.63" />
                    <SPLIT distance="400" swimtime="00:06:17.57" />
                    <SPLIT distance="500" swimtime="00:07:55.00" />
                    <SPLIT distance="600" swimtime="00:09:31.81" />
                    <SPLIT distance="700" swimtime="00:11:05.38" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="755" eventid="32" swimtime="00:01:14.39" lane="6" heatid="32002" />
                <RESULT resultid="756" eventid="34" swimtime="00:06:15.08" lane="4" heatid="34001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:22.62" />
                    <SPLIT distance="200" swimtime="00:03:01.60" />
                    <SPLIT distance="300" swimtime="00:04:39.27" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="200" birthdate="2004-01-01" gender="F" lastname="Placzek" firstname="Lilly" license="0">
              <RESULTS>
                <RESULT resultid="758" eventid="1" swimtime="00:00:19.90" lane="3" heatid="1015" />
                <RESULT resultid="763" eventid="5" swimtime="00:00:49.82" lane="4" heatid="5004" />
                <RESULT resultid="1409" eventid="7" swimtime="00:00:19.71" lane="7" heatid="7001" />
                <RESULT resultid="759" eventid="13" swimtime="00:00:41.28" lane="5" heatid="13007" />
                <RESULT resultid="760" eventid="19" swimtime="00:03:41.76" lane="5" heatid="19002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:50.99" />
                    <SPLIT distance="200" swimtime="00:01:47.62" />
                    <SPLIT distance="300" swimtime="00:02:46.74" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1497" eventid="21" swimtime="00:00:41.53" lane="2" heatid="21001" />
                <RESULT resultid="761" eventid="31" swimtime="00:00:45.24" lane="6" heatid="31016" />
                <RESULT resultid="762" eventid="37" swimtime="00:00:18.07" lane="5" heatid="37007" />
                <RESULT resultid="764" eventid="39" swimtime="00:00:22.72" lane="4" heatid="39004" />
                <RESULT resultid="1557" eventid="45" swimtime="00:00:17.78" lane="1" heatid="45001" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="201" birthdate="2002-01-01" gender="F" lastname="Klabunde" firstname="Lotte" license="0">
              <RESULTS>
                <RESULT resultid="765" eventid="1" swimtime="00:00:21.13" lane="2" heatid="1015" />
                <RESULT resultid="767" eventid="15" swimtime="00:01:42.35" lane="6" heatid="15011">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:50.23" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="768" eventid="27" swimtime="00:03:44.95" lane="8" heatid="27001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:51.96" />
                    <SPLIT distance="200" swimtime="00:01:49.22" />
                    <SPLIT distance="300" swimtime="00:02:48.75" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="769" eventid="31" swimtime="00:00:45.86" lane="6" heatid="31015" />
                <RESULT resultid="771" eventid="37" swimtime="00:00:19.05" lane="3" heatid="37005" />
                <RESULT resultid="770" eventid="43" swimtime="00:03:44.90" lane="8" heatid="43001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:53.40" />
                    <SPLIT distance="200" swimtime="00:01:50.21" />
                    <SPLIT distance="300" swimtime="00:02:48.43" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="202" birthdate="1986-01-01" gender="F" lastname="Klar" firstname="Margarethe" license="0">
              <RESULTS>
                <RESULT resultid="772" eventid="1" swimtime="00:00:28.12" lane="1" heatid="1006" />
                <RESULT resultid="773" eventid="13" swimtime="00:00:56.88" lane="2" heatid="13004" />
                <RESULT resultid="774" eventid="19" swimtime="00:04:28.51" lane="8" heatid="19002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:00.34" />
                    <SPLIT distance="200" swimtime="00:02:09.92" />
                    <SPLIT distance="300" swimtime="00:03:21.47" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="775" eventid="31" swimtime="00:01:00.99" lane="8" heatid="31007" />
                <RESULT resultid="776" eventid="33" swimtime="00:04:42.63" lane="1" heatid="33005">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:04.10" />
                    <SPLIT distance="200" swimtime="00:02:17.02" />
                    <SPLIT distance="300" swimtime="00:03:31.70" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="203" birthdate="2000-01-01" gender="F" lastname="Rütze" firstname="Michele" license="0">
              <RESULTS>
                <RESULT resultid="777" eventid="1" swimtime="00:00:19.59" lane="4" heatid="1015" />
                <RESULT resultid="1407" eventid="7" swimtime="00:00:18.65" lane="6" heatid="7001" />
                <RESULT resultid="778" eventid="13" swimtime="00:00:40.13" lane="4" heatid="13007" />
                <RESULT resultid="779" eventid="15" swimtime="00:01:36.13" lane="4" heatid="15012">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:45.95" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1494" eventid="21" swimtime="00:00:38.46" lane="5" heatid="21001" />
                <RESULT resultid="1515" eventid="23" swimtime="00:01:34.72" lane="5" heatid="23001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:46.18" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="780" eventid="31" swimtime="00:00:42.89" lane="4" heatid="31017" />
                <RESULT resultid="781" eventid="37" swimtime="00:00:17.28" lane="4" heatid="37008" />
                <RESULT resultid="1537" eventid="41" swimtime="00:00:40.95" lane="3" heatid="41001" />
                <RESULT resultid="1551" eventid="45" swimtime="00:00:17.18" lane="4" heatid="45001" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="204" birthdate="1978-01-01" gender="M" lastname="Hoffmann" firstname="Stefan" license="0">
              <RESULTS>
                <RESULT resultid="782" eventid="2" swimtime="00:00:22.61" lane="3" heatid="2007" />
                <RESULT resultid="785" eventid="6" swimtime="00:00:51.97" lane="7" heatid="6003" />
                <RESULT resultid="783" eventid="14" swimtime="00:00:46.54" lane="3" heatid="14003" />
                <RESULT resultid="784" eventid="38" swimtime="00:00:19.28" lane="1" heatid="38006" />
                <RESULT resultid="786" eventid="40" swimtime="00:00:24.11" lane="5" heatid="40003" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY number="3" gender="F" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="742" eventid="11" swimtime="00:06:44.78" lane="5" heatid="11003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:47.21" />
                    <SPLIT distance="200" swimtime="00:01:38.50" />
                    <SPLIT distance="300" swimtime="00:02:26.63" />
                    <SPLIT distance="400" swimtime="00:03:20.31" />
                    <SPLIT distance="500" swimtime="00:04:10.72" />
                    <SPLIT distance="600" swimtime="00:05:05.73" />
                    <SPLIT distance="700" swimtime="00:05:53.06" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="198" number="1" />
                    <RELAYPOSITION athleteid="201" number="2" />
                    <RELAYPOSITION athleteid="200" number="3" />
                    <RELAYPOSITION athleteid="203" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="3" gender="F" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="1383" eventid="48" swimtime="00:03:16.08" lane="5" heatid="48003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:45.40" />
                    <SPLIT distance="200" swimtime="00:01:31.60" />
                    <SPLIT distance="300" swimtime="00:02:33.49" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="200" number="1" />
                    <RELAYPOSITION athleteid="201" number="2" />
                    <RELAYPOSITION athleteid="202" number="3" />
                    <RELAYPOSITION athleteid="203" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB name="SG Finswimming Jena" nation="GER" region="35" code="174133">
          <ATHLETES>
            <ATHLETE athleteid="46" birthdate="2008-01-01" gender="M" lastname="Steininger" firstname="Bruno" license="0">
              <RESULTS>
                <RESULT resultid="135" eventid="14" swimtime="00:00:51.62" lane="3" heatid="14002" />
                <RESULT resultid="136" eventid="16" swimtime="00:01:55.40" lane="7" heatid="16005">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:56.47" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="137" eventid="20" swimtime="00:04:33.73" lane="6" heatid="20002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:02.24" />
                    <SPLIT distance="200" swimtime="00:02:13.31" />
                    <SPLIT distance="300" swimtime="00:03:25.65" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="138" eventid="34" swimtime="00:04:15.93" lane="8" heatid="34005">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:56.75" />
                    <SPLIT distance="200" swimtime="00:02:02.85" />
                    <SPLIT distance="300" swimtime="00:03:11.23" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="139" eventid="38" swimtime="00:00:20.63" lane="1" heatid="38004" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="47" birthdate="1999-01-01" gender="F" lastname="Jacke" firstname="Lena" license="0">
              <RESULTS>
                <RESULT resultid="140" eventid="3" swimtime="00:16:42.47" lane="3" heatid="3002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:01.80" />
                    <SPLIT distance="200" swimtime="00:02:05.66" />
                    <SPLIT distance="300" swimtime="00:03:13.30" />
                    <SPLIT distance="400" swimtime="00:04:18.49" />
                    <SPLIT distance="500" swimtime="00:05:28.07" />
                    <SPLIT distance="600" swimtime="00:06:34.24" />
                    <SPLIT distance="700" swimtime="00:07:44.41" />
                    <SPLIT distance="800" swimtime="00:08:50.92" />
                    <SPLIT distance="900" swimtime="00:10:01.04" />
                    <SPLIT distance="1000" swimtime="00:11:07.70" />
                    <SPLIT distance="1100" swimtime="00:12:17.87" />
                    <SPLIT distance="1200" swimtime="00:13:25.04" />
                    <SPLIT distance="1300" swimtime="00:14:34.95" />
                    <SPLIT distance="1400" swimtime="00:15:41.46" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="141" eventid="15" swimtime="00:01:54.57" lane="1" heatid="15009">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:55.61" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="142" eventid="17" swimtime="00:08:42.51" lane="6" heatid="17004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:01.74" />
                    <SPLIT distance="200" swimtime="00:02:05.75" />
                    <SPLIT distance="300" swimtime="00:03:13.84" />
                    <SPLIT distance="400" swimtime="00:04:18.91" />
                    <SPLIT distance="500" swimtime="00:05:28.70" />
                    <SPLIT distance="600" swimtime="00:06:33.83" />
                    <SPLIT distance="700" swimtime="00:07:41.91" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="143" eventid="31" swimtime="00:00:51.77" lane="7" heatid="31003" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="48" birthdate="2006-01-01" gender="F" lastname="Steininger" firstname="Liese" license="0">
              <RESULTS>
                <RESULT resultid="144" eventid="13" swimtime="00:00:57.69" lane="1" heatid="13002" />
                <RESULT resultid="145" eventid="19" swimtime="00:04:52.82" lane="8" heatid="19001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:06.04" />
                    <SPLIT distance="200" swimtime="00:02:20.84" />
                    <SPLIT distance="300" swimtime="00:03:37.41" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="146" eventid="31" swimtime="00:00:58.53" lane="5" heatid="31005" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="49" birthdate="2005-01-01" gender="F" lastname="Altenstein" firstname="Louise" license="0">
              <RESULTS>
                <RESULT resultid="147" eventid="3" swimtime="00:16:36.89" lane="4" heatid="3002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:57.03" />
                    <SPLIT distance="200" swimtime="00:01:59.91" />
                    <SPLIT distance="300" swimtime="00:03:05.59" />
                    <SPLIT distance="400" swimtime="00:04:08.30" />
                    <SPLIT distance="500" swimtime="00:05:16.28" />
                    <SPLIT distance="600" swimtime="00:06:21.48" />
                    <SPLIT distance="700" swimtime="00:07:30.87" />
                    <SPLIT distance="800" swimtime="00:08:37.83" />
                    <SPLIT distance="900" swimtime="00:09:48.28" />
                    <SPLIT distance="1000" swimtime="00:10:56.35" />
                    <SPLIT distance="1100" swimtime="00:12:06.21" />
                    <SPLIT distance="1200" swimtime="00:13:14.45" />
                    <SPLIT distance="1300" swimtime="00:14:26.38" />
                    <SPLIT distance="1400" swimtime="00:15:34.06" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="148" eventid="13" swimtime="00:00:47.51" lane="7" heatid="13006" />
                <RESULT resultid="149" eventid="17" swimtime="00:08:30.46" lane="2" heatid="17005">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:59.07" />
                    <SPLIT distance="200" swimtime="00:02:00.77" />
                    <SPLIT distance="300" swimtime="00:03:07.34" />
                    <SPLIT distance="400" swimtime="00:04:11.20" />
                    <SPLIT distance="500" swimtime="00:05:18.16" />
                    <SPLIT distance="600" swimtime="00:06:22.99" />
                    <SPLIT distance="700" swimtime="00:07:28.82" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="150" eventid="19" swimtime="00:04:03.93" lane="3" heatid="19002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:54.78" />
                    <SPLIT distance="200" swimtime="00:01:57.96" />
                    <SPLIT distance="300" swimtime="00:03:03.34" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="151" eventid="33" swimtime="00:04:00.64" lane="1" heatid="33007">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:55.01" />
                    <SPLIT distance="200" swimtime="00:01:55.11" />
                    <SPLIT distance="300" swimtime="00:02:59.22" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="152" eventid="37" swimtime="00:00:19.96" lane="8" heatid="37007" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="50" birthdate="2009-01-01" gender="F" lastname="Steininger" firstname="Magda" license="0">
              <RESULTS>
                <RESULT resultid="153" eventid="1" swimtime="00:00:24.94" lane="5" heatid="1008" />
                <RESULT resultid="154" eventid="13" swimtime="00:00:58.62" lane="7" heatid="13003" />
                <RESULT resultid="155" eventid="15" swimtime="00:02:10.50" lane="2" heatid="15005">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:03.00" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="156" eventid="31" swimtime="00:00:56.29" lane="1" heatid="31007" />
                <RESULT resultid="157" eventid="37" status="DNS" swimtime="00:00:00.00" lane="7" heatid="37002" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="51" birthdate="2005-01-01" gender="M" lastname="Preuß" firstname="Marek" license="0">
              <RESULTS>
                <RESULT resultid="158" eventid="10" swimtime="00:14:59.22" lane="6" heatid="10001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:56.86" />
                    <SPLIT distance="200" swimtime="00:01:57.12" />
                    <SPLIT distance="300" swimtime="00:02:59.04" />
                    <SPLIT distance="400" swimtime="00:03:56.90" />
                    <SPLIT distance="500" swimtime="00:04:59.14" />
                    <SPLIT distance="600" swimtime="00:05:59.21" />
                    <SPLIT distance="700" swimtime="00:07:02.79" />
                    <SPLIT distance="800" swimtime="00:07:59.82" />
                    <SPLIT distance="900" swimtime="00:09:04.42" />
                    <SPLIT distance="1000" swimtime="00:10:05.08" />
                    <SPLIT distance="1100" swimtime="00:11:01.96" />
                    <SPLIT distance="1200" swimtime="00:12:05.56" />
                    <SPLIT distance="1300" swimtime="00:13:07.33" />
                    <SPLIT distance="1400" swimtime="00:14:09.78" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="159" eventid="14" swimtime="00:00:43.96" lane="7" heatid="14005" />
                <RESULT resultid="160" eventid="28" swimtime="00:03:31.29" lane="6" heatid="28001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:49.76" />
                    <SPLIT distance="200" swimtime="00:01:42.74" />
                    <SPLIT distance="300" swimtime="00:02:37.14" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="161" eventid="34" swimtime="00:03:43.27" lane="5" heatid="34006">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:51.60" />
                    <SPLIT distance="200" swimtime="00:01:48.20" />
                    <SPLIT distance="300" swimtime="00:02:46.64" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="162" eventid="38" swimtime="00:00:19.24" lane="2" heatid="38006" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY number="1" gender="F" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="133" eventid="11" swimtime="00:08:04.05" lane="2" heatid="11002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:54.11" />
                    <SPLIT distance="200" swimtime="00:01:50.57" />
                    <SPLIT distance="300" swimtime="00:02:52.63" />
                    <SPLIT distance="400" swimtime="00:04:01.60" />
                    <SPLIT distance="500" swimtime="00:05:03.52" />
                    <SPLIT distance="600" swimtime="00:06:08.78" />
                    <SPLIT distance="700" swimtime="00:07:04.36" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="49" number="1" />
                    <RELAYPOSITION athleteid="50" number="2" />
                    <RELAYPOSITION athleteid="48" number="3" />
                    <RELAYPOSITION athleteid="47" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT resultid="134" eventid="48" swimtime="00:03:32.86" lane="7" heatid="48002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:48.47" />
                    <SPLIT distance="200" swimtime="00:01:44.44" />
                    <SPLIT distance="300" swimtime="00:02:41.78" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="49" number="1" />
                    <RELAYPOSITION athleteid="50" number="2" />
                    <RELAYPOSITION athleteid="48" number="3" />
                    <RELAYPOSITION athleteid="47" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB name="SSC Halle" nation="GER" region="27" code="0">
          <ATHLETES>
            <ATHLETE athleteid="284" birthdate="2007-01-01" gender="M" lastname="Koch" firstname="Elias" license="0">
              <RESULTS>
                <RESULT resultid="1081" eventid="2" swimtime="00:00:20.47" lane="1" heatid="2008" />
                <RESULT resultid="1082" eventid="14" swimtime="00:00:46.52" lane="2" heatid="14002" />
                <RESULT resultid="1083" eventid="32" swimtime="00:00:45.43" lane="5" heatid="32007" />
                <RESULT resultid="1084" eventid="38" swimtime="00:00:18.67" lane="3" heatid="38005" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="285" birthdate="2008-01-01" gender="M" lastname="Baumbach" firstname="Felix" license="0">
              <RESULTS>
                <RESULT resultid="1085" eventid="16" swimtime="00:01:54.60" lane="4" heatid="16005">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:55.06" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1086" eventid="18" swimtime="00:08:50.45" lane="4" heatid="18002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:02.28" />
                    <SPLIT distance="200" swimtime="00:02:09.15" />
                    <SPLIT distance="300" swimtime="00:03:17.05" />
                    <SPLIT distance="400" swimtime="00:04:25.85" />
                    <SPLIT distance="500" swimtime="00:05:34.14" />
                    <SPLIT distance="600" swimtime="00:06:42.59" />
                    <SPLIT distance="700" swimtime="00:07:48.77" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1087" eventid="32" swimtime="00:00:51.50" lane="2" heatid="32007" />
                <RESULT resultid="1088" eventid="34" swimtime="00:04:06.00" lane="4" heatid="34004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:57.76" />
                    <SPLIT distance="200" swimtime="00:02:01.86" />
                    <SPLIT distance="300" swimtime="00:03:06.18" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="286" birthdate="2011-01-01" gender="M" lastname="Reinicke" firstname="Jakob" license="0">
              <RESULTS>
                <RESULT resultid="1089" eventid="2" swimtime="00:00:25.91" lane="2" heatid="2002" />
                <RESULT resultid="1090" eventid="16" swimtime="00:02:11.62" lane="3" heatid="16003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:03.68" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1091" eventid="32" swimtime="00:01:00.47" lane="1" heatid="32003" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="287" birthdate="1984-01-01" gender="M" lastname="Hoffmann" firstname="Jörg" license="0">
              <RESULTS>
                <RESULT resultid="1092" eventid="2" swimtime="00:00:22.34" lane="2" heatid="2004" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="288" birthdate="2010-01-01" gender="M" lastname="Harms" firstname="Justus" license="0">
              <RESULTS>
                <RESULT resultid="1093" eventid="2" swimtime="00:00:27.63" lane="4" heatid="2002" />
                <RESULT resultid="1094" eventid="32" swimtime="00:01:01.79" lane="7" heatid="32003" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="289" birthdate="2007-01-01" gender="F" lastname="Gallitz" firstname="Laura" license="0">
              <RESULTS>
                <RESULT resultid="1095" eventid="1" swimtime="00:00:24.56" lane="2" heatid="1006" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="290" birthdate="2006-01-01" gender="F" lastname="Dietrich" firstname="Lea" license="0">
              <RESULTS>
                <RESULT resultid="1096" eventid="1" swimtime="00:00:20.58" lane="8" heatid="1015" />
                <RESULT resultid="1097" eventid="15" swimtime="00:01:49.17" lane="5" heatid="15008">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:52.34" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1098" eventid="31" swimtime="00:00:47.16" lane="7" heatid="31014" />
                <RESULT resultid="1099" eventid="37" swimtime="00:00:19.31" lane="7" heatid="37006" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="291" birthdate="2007-01-01" gender="F" lastname="Gerlach" firstname="Meret" license="0">
              <RESULTS>
                <RESULT resultid="1100" eventid="3" swimtime="00:16:40.49" lane="7" heatid="3002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:59.39" />
                    <SPLIT distance="200" swimtime="00:02:07.08" />
                    <SPLIT distance="300" swimtime="00:03:15.33" />
                    <SPLIT distance="400" swimtime="00:04:22.67" />
                    <SPLIT distance="500" swimtime="00:05:31.02" />
                    <SPLIT distance="600" swimtime="00:06:38.07" />
                    <SPLIT distance="700" swimtime="00:07:44.18" />
                    <SPLIT distance="800" swimtime="00:08:52.29" />
                    <SPLIT distance="900" swimtime="00:09:59.83" />
                    <SPLIT distance="1000" swimtime="00:11:07.38" />
                    <SPLIT distance="1100" swimtime="00:12:14.32" />
                    <SPLIT distance="1200" swimtime="00:13:23.36" />
                    <SPLIT distance="1300" swimtime="00:14:30.67" />
                    <SPLIT distance="1400" swimtime="00:15:37.36" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1101" eventid="15" swimtime="00:01:49.51" lane="3" heatid="15008">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:53.46" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1102" eventid="17" swimtime="00:08:21.97" lane="1" heatid="17005">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:58.51" />
                    <SPLIT distance="200" swimtime="00:02:01.80" />
                    <SPLIT distance="300" swimtime="00:03:06.14" />
                    <SPLIT distance="400" swimtime="00:04:10.86" />
                    <SPLIT distance="500" swimtime="00:05:15.76" />
                    <SPLIT distance="600" swimtime="00:06:20.51" />
                    <SPLIT distance="700" swimtime="00:07:24.00" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1103" eventid="31" swimtime="00:00:49.03" lane="1" heatid="31012" />
                <RESULT resultid="1104" eventid="33" swimtime="00:03:58.53" lane="6" heatid="33005">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:56.32" />
                    <SPLIT distance="200" swimtime="00:01:57.58" />
                    <SPLIT distance="300" swimtime="00:02:58.90" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="292" birthdate="2009-01-01" gender="M" lastname="Gaudig" firstname="Paul" license="0">
              <RESULTS>
                <RESULT resultid="1105" eventid="2" swimtime="00:00:22.48" lane="8" heatid="2006" />
                <RESULT resultid="1106" eventid="32" status="DSQ" swimtime="00:00:53.30" lane="8" heatid="32006" comment="Falscher Start." />
                <RESULT resultid="1107" eventid="38" swimtime="00:00:22.06" lane="4" heatid="38002" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="293" birthdate="2011-01-01" gender="M" lastname="Frenzel" firstname="Tim" license="0">
              <RESULTS>
                <RESULT resultid="1108" eventid="2" swimtime="00:00:32.96" lane="6" heatid="2001" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="294" birthdate="2010-01-01" gender="M" lastname="Eichberg" firstname="Eric" license="0" />
          </ATHLETES>
          <RELAYS>
            <RELAY number="1" gender="X" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="1079" eventid="30" swimtime="00:01:25.51" lane="3" heatid="30003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:42.01" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="284" number="1" />
                    <RELAYPOSITION athleteid="291" number="2" />
                    <RELAYPOSITION athleteid="285" number="3" />
                    <RELAYPOSITION athleteid="290" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" gender="M" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="1080" eventid="12" swimtime="00:09:57.86" lane="3" heatid="12001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:13.59" />
                    <SPLIT distance="200" swimtime="00:02:30.95" />
                    <SPLIT distance="300" swimtime="00:03:48.78" />
                    <SPLIT distance="400" swimtime="00:05:07.86" />
                    <SPLIT distance="500" swimtime="00:06:11.59" />
                    <SPLIT distance="600" swimtime="00:07:24.51" />
                    <SPLIT distance="700" swimtime="00:08:39.84" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="293" number="1" />
                    <RELAYPOSITION athleteid="294" number="2" />
                    <RELAYPOSITION athleteid="286" number="3" />
                    <RELAYPOSITION athleteid="288" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB name="SSV Freiburg" nation="GER" region="33" code="0">
          <ATHLETES>
            <ATHLETE athleteid="11" birthdate="1968-01-01" gender="M" lastname="Rolker" firstname="Bernd" license="100810">
              <RESULTS>
                <RESULT resultid="54" eventid="10" swimtime="00:17:11.52" lane="1" heatid="10001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:01.54" />
                    <SPLIT distance="200" swimtime="00:02:08.76" />
                    <SPLIT distance="300" swimtime="00:03:15.99" />
                    <SPLIT distance="400" swimtime="00:04:23.75" />
                    <SPLIT distance="500" swimtime="00:05:31.35" />
                    <SPLIT distance="600" swimtime="00:06:39.82" />
                    <SPLIT distance="700" swimtime="00:07:49.34" />
                    <SPLIT distance="800" swimtime="00:08:58.63" />
                    <SPLIT distance="900" swimtime="00:10:07.89" />
                    <SPLIT distance="1000" swimtime="00:11:18.48" />
                    <SPLIT distance="1100" swimtime="00:12:29.45" />
                    <SPLIT distance="1200" swimtime="00:13:41.32" />
                    <SPLIT distance="1300" swimtime="00:14:53.01" />
                    <SPLIT distance="1400" swimtime="00:16:03.46" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="55" eventid="14" swimtime="00:00:53.32" lane="1" heatid="14002" />
                <RESULT resultid="56" eventid="18" swimtime="00:09:04.20" lane="7" heatid="18003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:04.91" />
                    <SPLIT distance="200" swimtime="00:02:13.13" />
                    <SPLIT distance="300" swimtime="00:03:21.84" />
                    <SPLIT distance="400" swimtime="00:04:30.94" />
                    <SPLIT distance="500" swimtime="00:05:40.55" />
                    <SPLIT distance="600" swimtime="00:06:49.95" />
                    <SPLIT distance="700" swimtime="00:07:57.91" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="57" eventid="34" swimtime="00:04:33.80" lane="5" heatid="34005">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:02.83" />
                    <SPLIT distance="200" swimtime="00:02:10.40" />
                    <SPLIT distance="300" swimtime="00:03:21.92" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="58" eventid="38" swimtime="00:00:23.55" lane="4" heatid="38001" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="12" birthdate="1998-01-01" gender="F" lastname="Köhn" firstname="Johanna" license="100810">
              <RESULTS>
                <RESULT resultid="59" eventid="9" swimtime="00:15:22.37" lane="2" heatid="9001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:55.92" />
                    <SPLIT distance="200" swimtime="00:01:55.51" />
                    <SPLIT distance="300" swimtime="00:02:55.94" />
                    <SPLIT distance="400" swimtime="00:03:56.59" />
                    <SPLIT distance="500" swimtime="00:04:57.69" />
                    <SPLIT distance="600" swimtime="00:05:59.60" />
                    <SPLIT distance="700" swimtime="00:07:02.04" />
                    <SPLIT distance="800" swimtime="00:08:04.84" />
                    <SPLIT distance="900" swimtime="00:09:07.93" />
                    <SPLIT distance="1000" swimtime="00:10:10.83" />
                    <SPLIT distance="1100" swimtime="00:11:13.82" />
                    <SPLIT distance="1200" swimtime="00:12:17.12" />
                    <SPLIT distance="1300" swimtime="00:13:20.26" />
                    <SPLIT distance="1400" swimtime="00:14:22.35" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="60" eventid="15" swimtime="00:01:45.53" lane="2" heatid="15010">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:51.69" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="61" eventid="27" swimtime="00:03:49.03" lane="1" heatid="27001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:54.16" />
                    <SPLIT distance="200" swimtime="00:01:51.51" />
                    <SPLIT distance="300" swimtime="00:02:50.74" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="62" eventid="31" swimtime="00:00:47.99" lane="5" heatid="31014" />
                <RESULT resultid="63" eventid="33" swimtime="00:03:46.86" lane="5" heatid="33007">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:54.15" />
                    <SPLIT distance="200" swimtime="00:01:51.62" />
                    <SPLIT distance="300" swimtime="00:02:50.69" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="13" birthdate="1980-01-01" gender="M" lastname="Schmidt" firstname="Sascha" license="100810">
              <RESULTS>
                <RESULT resultid="1382" eventid="2" swimtime="00:00:20.67" lane="8" heatid="2001" />
                <RESULT resultid="64" eventid="14" swimtime="00:00:42.86" lane="1" heatid="14006" />
                <RESULT resultid="65" eventid="16" swimtime="00:01:46.57" lane="8" heatid="16008">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:50.19" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="66" eventid="18" swimtime="00:08:44.11" lane="5" heatid="18003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:59.72" />
                    <SPLIT distance="200" swimtime="00:02:02.92" />
                    <SPLIT distance="300" swimtime="00:03:07.73" />
                    <SPLIT distance="400" swimtime="00:04:13.46" />
                    <SPLIT distance="500" swimtime="00:05:20.26" />
                    <SPLIT distance="600" swimtime="00:06:28.14" />
                    <SPLIT distance="700" swimtime="00:07:36.62" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="67" eventid="28" swimtime="00:03:41.79" lane="2" heatid="28001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:48.44" />
                    <SPLIT distance="200" swimtime="00:01:43.59" />
                    <SPLIT distance="300" swimtime="00:02:41.17" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="68" eventid="32" swimtime="00:00:46.13" lane="1" heatid="32008" />
                <RESULT resultid="69" eventid="34" swimtime="00:04:06.42" lane="4" heatid="34005">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:56.50" />
                    <SPLIT distance="200" swimtime="00:01:58.34" />
                    <SPLIT distance="300" swimtime="00:03:02.33" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="70" eventid="38" swimtime="00:00:18.93" lane="3" heatid="38006" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="14" birthdate="2000-01-01" gender="F" lastname="Köhn" firstname="Theresa" license="100810">
              <RESULTS>
                <RESULT resultid="71" eventid="13" swimtime="00:00:44.30" lane="6" heatid="13006" />
                <RESULT resultid="1491" eventid="21" status="WDR" swimtime="00:00:00.00" lane="0" heatid="21000" />
                <RESULT resultid="72" eventid="27" swimtime="00:03:41.07" lane="6" heatid="27001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:50.84" />
                    <SPLIT distance="200" swimtime="00:01:45.95" />
                    <SPLIT distance="300" swimtime="00:02:43.96" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="73" eventid="31" swimtime="00:00:47.75" lane="2" heatid="31014" />
                <RESULT resultid="74" eventid="37" swimtime="00:00:19.77" lane="8" heatid="37008" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="Tauchclub Harz" nation="GER" region="27" code="164127">
          <ATHLETES>
            <ATHLETE athleteid="318" birthdate="2011-01-01" gender="M" lastname="Beier" firstname="Anton" license="0">
              <RESULTS>
                <RESULT resultid="1187" eventid="2" swimtime="00:00:28.42" lane="4" heatid="2001" />
                <RESULT resultid="1188" eventid="16" swimtime="00:02:24.69" lane="4" heatid="16001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:06.03" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1189" eventid="32" swimtime="00:01:02.99" lane="7" heatid="32002" />
                <RESULT resultid="1190" eventid="34" swimtime="00:04:51.83" lane="1" heatid="34002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:08.72" />
                    <SPLIT distance="200" swimtime="00:02:24.15" />
                    <SPLIT distance="300" swimtime="00:03:41.50" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="319" birthdate="2007-01-01" gender="F" lastname="Risse" firstname="Elisabeth" license="164127390">
              <RESULTS>
                <RESULT resultid="1191" eventid="1" swimtime="00:00:22.38" lane="4" heatid="1010" />
                <RESULT resultid="1192" eventid="17" swimtime="00:08:59.83" lane="2" heatid="17004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:58.59" />
                    <SPLIT distance="200" swimtime="00:02:05.06" />
                    <SPLIT distance="300" swimtime="00:03:13.80" />
                    <SPLIT distance="400" swimtime="00:04:23.37" />
                    <SPLIT distance="500" swimtime="00:05:33.35" />
                    <SPLIT distance="600" swimtime="00:06:43.70" />
                    <SPLIT distance="700" swimtime="00:07:52.33" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1193" eventid="31" swimtime="00:00:49.94" lane="8" heatid="31013" />
                <RESULT resultid="1194" eventid="33" swimtime="00:04:15.03" lane="7" heatid="33006">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:57.70" />
                    <SPLIT distance="200" swimtime="00:02:03.84" />
                    <SPLIT distance="300" swimtime="00:03:10.03" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1195" eventid="37" swimtime="00:00:21.08" lane="5" heatid="37003" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="320" birthdate="2008-01-01" gender="M" lastname="Härter" firstname="Fynn" license="164127389">
              <RESULTS>
                <RESULT resultid="1196" eventid="2" swimtime="00:00:22.09" lane="8" heatid="2008" />
                <RESULT resultid="1197" eventid="16" swimtime="00:01:49.64" lane="5" heatid="16005">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:51.17" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1198" eventid="32" swimtime="00:00:50.11" lane="6" heatid="32007" />
                <RESULT resultid="1199" eventid="34" swimtime="00:04:05.26" lane="8" heatid="34006">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:56.15" />
                    <SPLIT distance="200" swimtime="00:02:01.01" />
                    <SPLIT distance="300" swimtime="00:03:05.42" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1200" eventid="38" swimtime="00:00:19.93" lane="3" heatid="38004" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="321" birthdate="2004-01-01" gender="M" lastname="Hass" firstname="Jan Henrik" license="0">
              <RESULTS>
                <RESULT resultid="1201" eventid="2" swimtime="00:00:19.35" lane="3" heatid="2009" />
                <RESULT resultid="1202" eventid="16" swimtime="00:01:44.99" lane="6" heatid="16007">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:48.58" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1203" eventid="32" swimtime="00:00:43.10" lane="8" heatid="32010" />
                <RESULT resultid="1204" eventid="38" swimtime="00:00:17.70" lane="1" heatid="38008" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="322" birthdate="2009-01-01" gender="F" lastname="Zündel" firstname="Marlene" license="164127391">
              <RESULTS>
                <RESULT resultid="1205" eventid="1" swimtime="00:00:22.94" lane="8" heatid="1008" />
                <RESULT resultid="1206" eventid="15" swimtime="00:01:57.09" lane="8" heatid="15007">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:55.90" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1207" eventid="31" swimtime="00:00:51.44" lane="4" heatid="31010" />
                <RESULT resultid="1208" eventid="33" swimtime="00:04:31.07" lane="5" heatid="33004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:00.48" />
                    <SPLIT distance="200" swimtime="00:02:12.06" />
                    <SPLIT distance="300" swimtime="00:03:22.06" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1209" eventid="37" swimtime="00:00:22.46" lane="1" heatid="37002" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="323" birthdate="2008-01-01" gender="F" lastname="Weißenborn" firstname="Marnie" license="0">
              <RESULTS>
                <RESULT resultid="1210" eventid="1" swimtime="00:00:21.63" lane="1" heatid="1014" />
                <RESULT resultid="1214" eventid="5" swimtime="00:00:54.56" lane="3" heatid="5004" />
                <RESULT resultid="1211" eventid="15" swimtime="00:01:48.67" lane="1" heatid="15010">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:52.78" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1212" eventid="31" swimtime="00:00:47.25" lane="8" heatid="31015" />
                <RESULT resultid="1213" eventid="37" swimtime="00:00:20.58" lane="1" heatid="37008" />
                <RESULT resultid="1215" eventid="39" status="DSQ" swimtime="00:00:25.07" lane="5" heatid="39003" comment="Falscher Start." />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="324" birthdate="2009-01-01" gender="M" lastname="Schmidt" firstname="Matty" license="164127">
              <RESULTS>
                <RESULT resultid="1216" eventid="2" swimtime="00:00:24.87" lane="7" heatid="2004" />
                <RESULT resultid="1217" eventid="16" swimtime="00:02:00.82" lane="1" heatid="16004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:01.26" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1218" eventid="32" swimtime="00:00:55.10" lane="8" heatid="32004" />
                <RESULT resultid="1219" eventid="34" swimtime="00:04:23.53" lane="5" heatid="34003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:04.21" />
                    <SPLIT distance="200" swimtime="00:02:14.59" />
                    <SPLIT distance="300" swimtime="00:03:21.16" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="325" birthdate="2003-01-01" gender="M" lastname="Dalichow" firstname="Noah" license="0">
              <RESULTS>
                <RESULT resultid="1220" eventid="2" swimtime="00:00:19.15" lane="3" heatid="2010" />
                <RESULT resultid="1221" eventid="14" swimtime="00:00:39.52" lane="6" heatid="14006" />
                <RESULT resultid="1511" eventid="22" swimtime="00:00:39.98" lane="8" heatid="22001" />
                <RESULT resultid="1222" eventid="32" swimtime="00:00:44.66" lane="5" heatid="32009" />
                <RESULT resultid="1223" eventid="38" swimtime="00:00:17.57" lane="3" heatid="38007" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="326" birthdate="2007-01-01" gender="F" lastname="von Gynz Rekowski" firstname="Sophie" license="164127383">
              <RESULTS>
                <RESULT resultid="1224" eventid="1" swimtime="00:00:23.11" lane="6" heatid="1009" />
                <RESULT resultid="1225" eventid="15" swimtime="00:02:01.33" lane="7" heatid="15007">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:57.63" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1226" eventid="31" swimtime="00:00:53.78" lane="1" heatid="31010" />
                <RESULT resultid="1227" eventid="33" status="DNS" swimtime="00:00:00.00" lane="7" heatid="33004" />
                <RESULT resultid="1228" eventid="37" swimtime="00:00:21.31" lane="1" heatid="37004" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY number="1" gender="F" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="1183" eventid="11" status="DSQ" swimtime="00:07:52.18" lane="4" heatid="11002" comment="Die 4. Sportlerin behinderte einen anderen Sportler auf Bahn 3.">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:54.40" />
                    <SPLIT distance="200" swimtime="00:01:50.69" />
                    <SPLIT distance="300" swimtime="00:02:47.40" />
                    <SPLIT distance="400" swimtime="00:03:51.85" />
                    <SPLIT distance="500" swimtime="00:04:51.03" />
                    <SPLIT distance="600" swimtime="00:05:54.48" />
                    <SPLIT distance="700" swimtime="00:06:47.98" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="323" number="1" />
                    <RELAYPOSITION athleteid="322" number="2" />
                    <RELAYPOSITION athleteid="326" number="3" />
                    <RELAYPOSITION athleteid="319" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT resultid="1184" eventid="48" swimtime="00:03:22.78" lane="8" heatid="48003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:48.00" />
                    <SPLIT distance="200" swimtime="00:01:40.21" />
                    <SPLIT distance="300" swimtime="00:02:32.46" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="323" number="1" />
                    <RELAYPOSITION athleteid="322" number="2" />
                    <RELAYPOSITION athleteid="326" number="3" />
                    <RELAYPOSITION athleteid="319" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="2" gender="X" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="1185" eventid="30" swimtime="00:01:29.18" lane="4" heatid="30003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:44.77" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="323" number="1" />
                    <RELAYPOSITION athleteid="324" number="2" />
                    <RELAYPOSITION athleteid="322" number="3" />
                    <RELAYPOSITION athleteid="320" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="3" gender="X" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="1186" eventid="30" swimtime="00:01:22.95" lane="7" heatid="30003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:40.93" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="325" number="1" />
                    <RELAYPOSITION athleteid="319" number="2" />
                    <RELAYPOSITION athleteid="326" number="3" />
                    <RELAYPOSITION athleteid="321" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB name="Tauchclub Heilbronn" nation="GER" region="32" code="124012">
          <ATHLETES>
            <ATHLETE athleteid="77" birthdate="2004-01-01" gender="F" lastname="Phillipp" firstname="Beeke Alea" license="0">
              <RESULTS>
                <RESULT resultid="255" eventid="1" swimtime="00:00:21.23" lane="5" heatid="1012" />
                <RESULT resultid="256" eventid="13" swimtime="00:00:45.89" lane="2" heatid="13007" />
                <RESULT resultid="257" eventid="15" swimtime="00:01:49.26" lane="7" heatid="15009">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:51.78" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="258" eventid="19" swimtime="00:04:09.11" lane="4" heatid="19001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:52.98" />
                    <SPLIT distance="200" swimtime="00:01:55.69" />
                    <SPLIT distance="300" swimtime="00:03:03.85" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="259" eventid="31" swimtime="00:00:47.45" lane="1" heatid="31014" />
                <RESULT resultid="260" eventid="37" swimtime="00:00:19.96" lane="4" heatid="37005" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="78" birthdate="2007-01-01" gender="M" lastname="Bilicz" firstname="Benedikt" license="0">
              <RESULTS>
                <RESULT resultid="261" eventid="2" swimtime="00:00:19.76" lane="3" heatid="2008" />
                <RESULT resultid="262" eventid="14" swimtime="00:00:45.02" lane="6" heatid="14003" />
                <RESULT resultid="263" eventid="16" swimtime="00:01:45.07" lane="1" heatid="16006">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:49.22" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="264" eventid="32" swimtime="00:00:45.50" lane="6" heatid="32008" />
                <RESULT resultid="265" eventid="38" swimtime="00:00:17.22" lane="5" heatid="38006" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="79" birthdate="2011-01-01" gender="M" lastname="Korb" firstname="Elias" license="0">
              <RESULTS>
                <RESULT resultid="266" eventid="2" swimtime="00:00:25.89" lane="6" heatid="2003" />
                <RESULT resultid="267" eventid="14" swimtime="00:00:51.85" lane="5" heatid="14001" />
                <RESULT resultid="268" eventid="16" swimtime="00:02:01.90" lane="5" heatid="16004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:00.29" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="269" eventid="20" swimtime="00:04:26.11" lane="2" heatid="20001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:03.37" />
                    <SPLIT distance="200" swimtime="00:02:12.84" />
                    <SPLIT distance="300" swimtime="00:03:22.48" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="270" eventid="32" swimtime="00:00:56.77" lane="6" heatid="32004" />
                <RESULT resultid="271" eventid="34" swimtime="00:04:14.93" lane="5" heatid="34004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:01.03" />
                    <SPLIT distance="200" swimtime="00:02:07.21" />
                    <SPLIT distance="300" swimtime="00:03:13.13" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="272" eventid="36" swimtime="00:00:24.21" lane="5" heatid="36001" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="80" birthdate="2009-01-01" gender="F" lastname="Hölzer" firstname="Elisa" license="0">
              <RESULTS>
                <RESULT resultid="273" eventid="1" swimtime="00:00:23.58" lane="1" heatid="1010" />
                <RESULT resultid="274" eventid="13" swimtime="00:00:53.29" lane="8" heatid="13004" />
                <RESULT resultid="275" eventid="15" swimtime="00:01:59.36" lane="8" heatid="15008">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:55.89" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="276" eventid="19" swimtime="00:04:24.41" lane="2" heatid="19001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:59.13" />
                    <SPLIT distance="200" swimtime="00:02:08.50" />
                    <SPLIT distance="300" swimtime="00:03:19.15" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="277" eventid="31" swimtime="00:00:51.34" lane="7" heatid="31010" />
                <RESULT resultid="278" eventid="33" swimtime="00:04:18.44" lane="2" heatid="33005">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:58.88" />
                    <SPLIT distance="200" swimtime="00:02:06.07" />
                    <SPLIT distance="300" swimtime="00:03:13.59" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="279" eventid="37" swimtime="00:00:22.08" lane="6" heatid="37003" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="81" birthdate="2008-01-01" gender="F" lastname="Seidel" firstname="Esther-Sophie" license="0">
              <RESULTS>
                <RESULT resultid="280" eventid="1" swimtime="00:00:21.95" lane="6" heatid="1011" />
                <RESULT resultid="281" eventid="15" swimtime="00:01:58.57" lane="8" heatid="15006">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:56.09" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="282" eventid="31" swimtime="00:00:50.58" lane="3" heatid="31010" />
                <RESULT resultid="283" eventid="37" swimtime="00:00:20.90" lane="6" heatid="37004" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="82" birthdate="2008-01-01" gender="F" lastname="Grimm" firstname="Hannah" license="0">
              <RESULTS>
                <RESULT resultid="284" eventid="1" swimtime="00:00:23.81" lane="4" heatid="1008" />
                <RESULT resultid="285" eventid="13" swimtime="00:00:56.63" lane="8" heatid="13003" />
                <RESULT resultid="286" eventid="31" swimtime="00:00:54.32" lane="7" heatid="31007" />
                <RESULT resultid="287" eventid="37" status="DNS" swimtime="00:00:00.00" lane="6" heatid="37002" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="83" birthdate="2000-01-01" gender="F" lastname="Baier" firstname="Jessika" license="0">
              <RESULTS>
                <RESULT resultid="288" eventid="1" swimtime="00:00:22.90" lane="2" heatid="1009" />
                <RESULT resultid="289" eventid="13" swimtime="00:00:51.63" lane="5" heatid="13004" />
                <RESULT resultid="290" eventid="15" swimtime="00:02:04.26" lane="4" heatid="15006">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:56.50" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="291" eventid="31" swimtime="00:00:52.04" lane="1" heatid="31009" />
                <RESULT resultid="292" eventid="37" swimtime="00:00:21.26" lane="3" heatid="37003" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="84" birthdate="2004-01-01" gender="F" lastname="Ruedel" firstname="Leona" license="0">
              <RESULTS>
                <RESULT resultid="293" eventid="1" swimtime="00:00:21.73" lane="2" heatid="1012" />
                <RESULT resultid="294" eventid="13" swimtime="00:00:45.85" lane="2" heatid="13006" />
                <RESULT resultid="295" eventid="15" swimtime="00:01:47.54" lane="8" heatid="15011">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:52.35" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="296" eventid="31" swimtime="00:00:46.67" lane="2" heatid="31012" />
                <RESULT resultid="297" eventid="37" swimtime="00:00:19.14" lane="7" heatid="37007" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="85" birthdate="2004-01-01" gender="M" lastname="Rist" firstname="Marc" license="0">
              <RESULTS>
                <RESULT resultid="298" eventid="2" swimtime="00:00:21.98" lane="5" heatid="2007" />
                <RESULT resultid="299" eventid="16" swimtime="00:01:50.01" lane="8" heatid="16006">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:53.76" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="300" eventid="18" swimtime="00:08:36.07" lane="8" heatid="18003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:59.48" />
                    <SPLIT distance="200" swimtime="00:02:04.41" />
                    <SPLIT distance="300" swimtime="00:03:10.86" />
                    <SPLIT distance="400" swimtime="00:04:17.57" />
                    <SPLIT distance="500" swimtime="00:05:24.33" />
                    <SPLIT distance="600" swimtime="00:06:30.66" />
                    <SPLIT distance="700" swimtime="00:07:36.06" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="301" eventid="32" swimtime="00:00:48.69" lane="6" heatid="32006" />
                <RESULT resultid="302" eventid="34" swimtime="00:04:09.54" lane="1" heatid="34006">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:56.13" />
                    <SPLIT distance="200" swimtime="00:02:01.91" />
                    <SPLIT distance="300" swimtime="00:03:08.35" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="86" birthdate="2011-01-01" gender="F" lastname="Jung" firstname="Sarah" license="0">
              <RESULTS>
                <RESULT resultid="303" eventid="1" swimtime="00:00:28.24" lane="8" heatid="1002" />
                <RESULT resultid="304" eventid="15" swimtime="00:02:28.39" lane="1" heatid="15002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:14.07" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="305" eventid="31" swimtime="00:01:04.93" lane="6" heatid="31002" />
                <RESULT resultid="306" eventid="35" swimtime="00:00:28.72" lane="2" heatid="35001" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="87" birthdate="2002-01-01" gender="M" lastname="Bauer" firstname="Sebastian" license="0">
              <RESULTS>
                <RESULT resultid="307" eventid="2" swimtime="00:00:23.52" lane="5" heatid="2006" />
                <RESULT resultid="308" eventid="18" swimtime="00:08:45.59" lane="1" heatid="18003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:59.77" />
                    <SPLIT distance="200" swimtime="00:02:05.23" />
                    <SPLIT distance="300" swimtime="00:03:11.37" />
                    <SPLIT distance="400" swimtime="00:04:17.81" />
                    <SPLIT distance="500" swimtime="00:05:25.22" />
                    <SPLIT distance="600" swimtime="00:06:33.09" />
                    <SPLIT distance="700" swimtime="00:07:40.75" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="309" eventid="32" swimtime="00:00:52.53" lane="5" heatid="32006" />
                <RESULT resultid="310" eventid="34" swimtime="00:04:12.81" lane="2" heatid="34005">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:58.09" />
                    <SPLIT distance="200" swimtime="00:02:02.14" />
                    <SPLIT distance="300" swimtime="00:03:07.90" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="88" birthdate="2009-01-01" gender="F" lastname="Rettig" firstname="Sina" license="0">
              <RESULTS>
                <RESULT resultid="311" eventid="1" swimtime="00:00:24.69" lane="4" heatid="1006" />
                <RESULT resultid="312" eventid="13" swimtime="00:01:02.98" lane="4" heatid="13001" />
                <RESULT resultid="313" eventid="15" swimtime="00:02:10.99" lane="4" heatid="15003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:02.81" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="314" eventid="31" swimtime="00:00:56.78" lane="3" heatid="31006" />
                <RESULT resultid="315" eventid="37" swimtime="00:00:23.77" lane="4" heatid="37001" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="89" birthdate="2003-01-01" gender="M" lastname="Fabriz" firstname="Tobias" license="0">
              <RESULTS>
                <RESULT resultid="316" eventid="2" swimtime="00:00:19.66" lane="7" heatid="2010" />
                <RESULT resultid="317" eventid="14" swimtime="00:00:41.77" lane="2" heatid="14005" />
                <RESULT resultid="318" eventid="32" swimtime="00:00:43.63" lane="3" heatid="32009" />
                <RESULT resultid="319" eventid="38" swimtime="00:00:17.05" lane="6" heatid="38007" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY number="1" gender="F" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="249" eventid="11" swimtime="00:08:15.07" lane="6" heatid="11002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:59.99" />
                    <SPLIT distance="200" swimtime="00:02:09.53" />
                    <SPLIT distance="300" swimtime="00:03:10.34" />
                    <SPLIT distance="400" swimtime="00:04:18.06" />
                    <SPLIT distance="500" swimtime="00:05:12.15" />
                    <SPLIT distance="600" swimtime="00:06:15.53" />
                    <SPLIT distance="700" swimtime="00:07:11.24" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="88" number="1" />
                    <RELAYPOSITION athleteid="82" number="2" />
                    <RELAYPOSITION athleteid="81" number="3" />
                    <RELAYPOSITION athleteid="80" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT resultid="250" eventid="48" swimtime="00:03:31.99" lane="6" heatid="48002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:56.09" />
                    <SPLIT distance="200" swimtime="00:01:49.84" />
                    <SPLIT distance="300" swimtime="00:02:40.24" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="88" number="1" />
                    <RELAYPOSITION athleteid="82" number="2" />
                    <RELAYPOSITION athleteid="81" number="3" />
                    <RELAYPOSITION athleteid="80" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="2" gender="M" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="251" eventid="12" swimtime="00:07:40.91" lane="2" heatid="12002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:56.14" />
                    <SPLIT distance="200" swimtime="00:01:58.41" />
                    <SPLIT distance="300" swimtime="00:02:51.85" />
                    <SPLIT distance="400" swimtime="00:03:49.16" />
                    <SPLIT distance="500" swimtime="00:04:49.48" />
                    <SPLIT distance="600" swimtime="00:05:54.23" />
                    <SPLIT distance="700" swimtime="00:06:43.07" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="87" number="1" />
                    <RELAYPOSITION athleteid="85" number="2" />
                    <RELAYPOSITION athleteid="79" number="3" />
                    <RELAYPOSITION athleteid="78" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="3" gender="X" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="252" eventid="30" swimtime="00:01:21.91" lane="5" heatid="30003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:40.36" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="89" number="1" />
                    <RELAYPOSITION athleteid="85" number="2" />
                    <RELAYPOSITION athleteid="84" number="3" />
                    <RELAYPOSITION athleteid="77" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="4" gender="X" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="253" eventid="30" swimtime="00:01:28.79" lane="1" heatid="30003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:47.38" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="81" number="1" />
                    <RELAYPOSITION athleteid="79" number="2" />
                    <RELAYPOSITION athleteid="80" number="3" />
                    <RELAYPOSITION athleteid="78" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="5" gender="M" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="254" eventid="49" swimtime="00:03:12.61" lane="7" heatid="49002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:55.79" />
                    <SPLIT distance="200" swimtime="00:01:44.94" />
                    <SPLIT distance="300" swimtime="00:02:29.61" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="79" number="1" />
                    <RELAYPOSITION athleteid="85" number="2" />
                    <RELAYPOSITION athleteid="78" number="3" />
                    <RELAYPOSITION athleteid="89" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB name="Tauchclub NEMO Plauen e.V." nation="GER" region="20" code="0">
          <ATHLETES>
            <ATHLETE athleteid="271" birthdate="2009-01-01" gender="F" lastname="Troppschuh" firstname="Hannah" license="0">
              <RESULTS>
                <RESULT resultid="1028" eventid="1" swimtime="00:00:21.19" lane="1" heatid="1013" />
                <RESULT resultid="1029" eventid="13" swimtime="00:00:44.57" lane="6" heatid="13007" />
                <RESULT resultid="1500" eventid="21" swimtime="00:00:43.91" lane="8" heatid="21001" />
                <RESULT resultid="1030" eventid="27" swimtime="00:03:40.88" lane="7" heatid="27001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:50.96" />
                    <SPLIT distance="200" swimtime="00:01:47.26" />
                    <SPLIT distance="300" swimtime="00:02:46.87" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1031" eventid="31" swimtime="00:00:47.44" lane="1" heatid="31017" />
                <RESULT resultid="1032" eventid="37" swimtime="00:00:19.04" lane="2" heatid="37008" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="272" birthdate="2003-01-01" gender="F" lastname="Prochaska" firstname="Julia" license="0">
              <RESULTS>
                <RESULT resultid="1033" eventid="1" swimtime="00:00:22.95" lane="2" heatid="1011" />
                <RESULT resultid="1034" eventid="13" swimtime="00:00:48.62" lane="7" heatid="13005" />
                <RESULT resultid="1035" eventid="31" swimtime="00:00:51.79" lane="7" heatid="31011" />
                <RESULT resultid="1036" eventid="37" swimtime="00:00:20.60" lane="7" heatid="37005" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="273" birthdate="1972-01-01" gender="M" lastname="Gräf" firstname="Sven" license="0">
              <RESULTS>
                <RESULT resultid="1037" eventid="2" status="DNS" swimtime="00:00:00.00" lane="6" heatid="2008" />
                <RESULT resultid="1038" eventid="6" status="DNS" swimtime="00:00:00.00" lane="4" heatid="6004" />
                <RESULT resultid="1039" eventid="40" status="DNS" swimtime="00:00:00.00" lane="8" heatid="40004" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="Tauchclub Oberspree e.V." nation="GER" region="21" code="3410800">
          <ATHLETES>
            <ATHLETE athleteid="67" birthdate="2009-01-01" gender="F" lastname="Kießling" firstname="Romy" license="0">
              <RESULTS>
                <RESULT resultid="222" eventid="1" swimtime="00:00:28.41" lane="8" heatid="1005" />
                <RESULT resultid="223" eventid="13" swimtime="00:00:57.81" lane="6" heatid="13002" />
                <RESULT resultid="224" eventid="15" swimtime="00:02:18.83" lane="8" heatid="15004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:06.01" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="225" eventid="17" status="DSQ" swimtime="00:00:00.00" lane="2" heatid="17002" comment="Aufgegeben nach 400 Meter.">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:08.68" />
                    <SPLIT distance="200" swimtime="00:02:25.23" />
                    <SPLIT distance="300" swimtime="00:03:43.75" />
                    <SPLIT distance="400" swimtime="00:05:05.38" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="226" eventid="31" swimtime="00:01:02.09" lane="4" heatid="31004" />
                <RESULT resultid="227" eventid="33" swimtime="00:04:50.92" lane="2" heatid="33002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:08.17" />
                    <SPLIT distance="200" swimtime="00:02:23.10" />
                    <SPLIT distance="300" swimtime="00:03:39.53" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="Tauchclub Potsdam" nation="GER" region="19" code="134111">
          <ATHLETES>
            <ATHLETE athleteid="15" birthdate="2003-01-01" gender="F" lastname="Junghans" firstname="Chiara" license="0">
              <RESULTS>
                <RESULT resultid="75" eventid="1" swimtime="00:00:21.47" lane="6" heatid="1012" />
                <RESULT resultid="80" eventid="5" swimtime="00:00:54.47" lane="7" heatid="5004" />
                <RESULT resultid="76" eventid="15" swimtime="00:01:42.74" lane="2" heatid="15011">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:49.09" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="77" eventid="25" swimtime="00:08:07.34" lane="8" heatid="25001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:55.37" />
                    <SPLIT distance="200" swimtime="00:01:55.33" />
                    <SPLIT distance="300" swimtime="00:02:56.82" />
                    <SPLIT distance="400" swimtime="00:03:58.84" />
                    <SPLIT distance="500" swimtime="00:05:01.59" />
                    <SPLIT distance="600" swimtime="00:06:04.21" />
                    <SPLIT distance="700" swimtime="00:07:06.87" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="78" eventid="31" swimtime="00:00:46.09" lane="8" heatid="31017" />
                <RESULT resultid="79" eventid="33" swimtime="00:03:48.04" lane="3" heatid="33007">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:53.25" />
                    <SPLIT distance="200" swimtime="00:01:50.88" />
                    <SPLIT distance="300" swimtime="00:02:50.28" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="81" eventid="39" swimtime="00:00:25.27" lane="8" heatid="39004" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="16" birthdate="1997-01-01" gender="F" lastname="Starke" firstname="Juliane" license="0">
              <RESULTS>
                <RESULT resultid="82" eventid="1" swimtime="00:00:21.68" lane="8" heatid="1012" />
                <RESULT resultid="87" eventid="5" swimtime="00:00:54.07" lane="2" heatid="5004" />
                <RESULT resultid="83" eventid="15" swimtime="00:01:42.30" lane="8" heatid="15012">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:49.29" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="84" eventid="19" swimtime="00:03:52.56" lane="7" heatid="19002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:53.35" />
                    <SPLIT distance="200" swimtime="00:01:53.40" />
                    <SPLIT distance="300" swimtime="00:02:54.28" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="85" eventid="31" swimtime="00:00:46.50" lane="6" heatid="31014" />
                <RESULT resultid="86" eventid="33" swimtime="00:03:46.03" lane="6" heatid="33007">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:53.26" />
                    <SPLIT distance="200" swimtime="00:01:51.35" />
                    <SPLIT distance="300" swimtime="00:02:50.07" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="88" eventid="39" swimtime="00:00:24.93" lane="7" heatid="39004" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="Tauchsport Döbeln" nation="GER" region="20" code="154104000">
          <ATHLETES>
            <ATHLETE athleteid="59" birthdate="2006-01-01" gender="M" lastname="Noack" firstname="Christopher" license="0">
              <RESULTS>
                <RESULT resultid="174" eventid="2" status="DNS" swimtime="00:00:00.00" lane="3" heatid="2005" />
                <RESULT resultid="177" eventid="6" status="DNS" swimtime="00:00:00.00" lane="7" heatid="6002" />
                <RESULT resultid="175" eventid="32" status="DNS" swimtime="00:00:00.00" lane="1" heatid="32005" />
                <RESULT resultid="176" eventid="38" status="DNS" swimtime="00:00:00.00" lane="3" heatid="38002" />
                <RESULT resultid="178" eventid="40" status="DNS" swimtime="00:00:00.00" lane="4" heatid="40002" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="60" birthdate="1973-01-01" gender="M" lastname="Winkler" firstname="Daniel" license="0">
              <RESULTS>
                <RESULT resultid="179" eventid="2" swimtime="00:00:23.27" lane="1" heatid="2006" />
                <RESULT resultid="185" eventid="6" swimtime="00:00:58.60" lane="3" heatid="6002" />
                <RESULT resultid="180" eventid="14" swimtime="00:00:47.65" lane="4" heatid="14002" />
                <RESULT resultid="181" eventid="16" swimtime="00:01:58.34" lane="3" heatid="16004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:55.45" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="182" eventid="20" swimtime="00:04:24.10" lane="8" heatid="20002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:59.35" />
                    <SPLIT distance="200" swimtime="00:02:11.17" />
                    <SPLIT distance="300" swimtime="00:03:21.29" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="183" eventid="32" swimtime="00:00:50.92" lane="6" heatid="32005" />
                <RESULT resultid="184" eventid="38" swimtime="00:00:20.33" lane="4" heatid="38003" />
                <RESULT resultid="186" eventid="40" swimtime="00:00:25.22" lane="5" heatid="40002" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="61" birthdate="2003-01-01" gender="M" lastname="Elenkow" firstname="Felix" license="0">
              <RESULTS>
                <RESULT resultid="187" eventid="2" swimtime="00:00:20.14" lane="2" heatid="2009" />
                <RESULT resultid="190" eventid="6" swimtime="00:00:51.40" lane="6" heatid="6004" />
                <RESULT resultid="188" eventid="32" swimtime="00:00:44.64" lane="1" heatid="32010" />
                <RESULT resultid="189" eventid="38" swimtime="00:00:18.87" lane="6" heatid="38002" />
                <RESULT resultid="191" eventid="40" swimtime="00:00:23.11" lane="5" heatid="40004" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="62" birthdate="1956-01-01" gender="M" lastname="Mönch" firstname="Helmut" license="0">
              <RESULTS>
                <RESULT resultid="192" eventid="2" swimtime="00:00:25.69" lane="7" heatid="2001" />
                <RESULT resultid="193" eventid="14" swimtime="00:00:53.73" lane="1" heatid="14001" />
                <RESULT resultid="194" eventid="20" swimtime="00:04:47.46" lane="5" heatid="20001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:03.70" />
                    <SPLIT distance="200" swimtime="00:02:17.87" />
                    <SPLIT distance="300" swimtime="00:03:33.69" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="195" eventid="32" swimtime="00:00:58.09" lane="3" heatid="32001" />
                <RESULT resultid="196" eventid="38" swimtime="00:00:23.10" lane="6" heatid="38001" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="63" birthdate="1962-01-01" gender="M" lastname="Muth" firstname="Henrik" license="0">
              <RESULTS>
                <RESULT resultid="197" eventid="2" swimtime="00:00:23.53" lane="6" heatid="2006" />
                <RESULT resultid="198" eventid="4" status="DNS" swimtime="00:00:00.00" lane="2" heatid="4001" />
                <RESULT resultid="206" eventid="6" swimtime="00:00:58.24" lane="6" heatid="6001" />
                <RESULT resultid="199" eventid="14" swimtime="00:00:48.55" lane="7" heatid="14003" />
                <RESULT resultid="200" eventid="16" swimtime="00:02:01.07" lane="6" heatid="16003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:59.27" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="201" eventid="18" swimtime="00:09:30.07" lane="4" heatid="18001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:01.21" />
                    <SPLIT distance="200" swimtime="00:02:12.68" />
                    <SPLIT distance="300" swimtime="00:03:26.18" />
                    <SPLIT distance="400" swimtime="00:04:39.78" />
                    <SPLIT distance="500" swimtime="00:05:53.65" />
                    <SPLIT distance="600" swimtime="00:07:07.22" />
                    <SPLIT distance="700" swimtime="00:08:21.21" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="202" eventid="20" swimtime="00:04:14.18" lane="1" heatid="20002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:54.81" />
                    <SPLIT distance="200" swimtime="00:02:00.50" />
                    <SPLIT distance="300" swimtime="00:03:08.50" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="203" eventid="32" swimtime="00:00:52.75" lane="7" heatid="32006" />
                <RESULT resultid="204" eventid="34" status="DNF" swimtime="00:00:00.00" lane="7" heatid="34002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:01.98" />
                    <SPLIT distance="200" swimtime="00:02:12.74" />
                    <SPLIT distance="300" swimtime="00:03:42.20" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="205" eventid="38" status="DNS" swimtime="00:00:00.00" lane="6" heatid="38004" />
                <RESULT resultid="207" eventid="40" status="DNS" swimtime="00:00:00.00" lane="2" heatid="40001" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="Tauchsportclub Erfurt e.V." nation="GER" region="35" code="0">
          <ATHLETES>
            <ATHLETE athleteid="156" birthdate="2010-01-01" gender="F" lastname="Abe" firstname="Adina" license="0">
              <RESULTS>
                <RESULT resultid="570" eventid="1" swimtime="00:00:23.03" lane="4" heatid="1009" />
                <RESULT resultid="571" eventid="13" swimtime="00:00:50.40" lane="8" heatid="13007" />
                <RESULT resultid="572" eventid="15" swimtime="00:01:53.04" lane="6" heatid="15008">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:54.48" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="573" eventid="31" swimtime="00:00:50.42" lane="6" heatid="31011" />
                <RESULT resultid="574" eventid="35" swimtime="00:00:23.17" lane="5" heatid="35002" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="157" birthdate="2009-01-01" gender="F" lastname="Darzhaniia" firstname="Alisa" license="0">
              <RESULTS>
                <RESULT resultid="575" eventid="1" swimtime="00:00:22.56" lane="3" heatid="1012" />
                <RESULT resultid="581" eventid="5" swimtime="00:00:57.12" lane="1" heatid="5004" />
                <RESULT resultid="576" eventid="15" swimtime="00:01:52.04" lane="3" heatid="15009">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:53.67" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="577" eventid="17" swimtime="00:08:32.37" lane="7" heatid="17005">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:58.09" />
                    <SPLIT distance="200" swimtime="00:02:02.53" />
                    <SPLIT distance="300" swimtime="00:03:07.81" />
                    <SPLIT distance="400" swimtime="00:04:14.51" />
                    <SPLIT distance="500" swimtime="00:05:21.00" />
                    <SPLIT distance="600" swimtime="00:06:27.86" />
                    <SPLIT distance="700" swimtime="00:07:32.29" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="579" eventid="33" swimtime="00:04:01.80" lane="6" heatid="33006">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:54.76" />
                    <SPLIT distance="200" swimtime="00:01:58.03" />
                    <SPLIT distance="300" swimtime="00:03:02.25" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="580" eventid="37" swimtime="00:00:20.65" lane="5" heatid="37005" />
                <RESULT resultid="582" eventid="39" swimtime="00:00:26.18" lane="4" heatid="39003" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="158" birthdate="2004-01-01" gender="F" lastname="Möller" firstname="Amelie" license="0">
              <RESULTS>
                <RESULT resultid="583" eventid="5" swimtime="00:01:03.03" lane="5" heatid="5002" />
                <RESULT resultid="584" eventid="39" swimtime="00:00:28.89" lane="6" heatid="39002" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="159" birthdate="2009-01-01" gender="F" lastname="Zitzmann" firstname="Annalena" license="0">
              <RESULTS>
                <RESULT resultid="585" eventid="1" swimtime="00:00:22.46" lane="5" heatid="1010" />
                <RESULT resultid="586" eventid="13" swimtime="00:00:50.73" lane="6" heatid="13004" />
                <RESULT resultid="587" eventid="15" swimtime="00:01:58.13" lane="5" heatid="15006">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:57.73" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="588" eventid="31" swimtime="00:00:50.81" lane="1" heatid="31011" />
                <RESULT resultid="589" eventid="37" swimtime="00:00:21.79" lane="2" heatid="37002" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="160" birthdate="2010-01-01" gender="M" lastname="Blumenstein" firstname="Einar" license="0">
              <RESULTS>
                <RESULT resultid="590" eventid="2" swimtime="00:00:26.68" lane="8" heatid="2002" />
                <RESULT resultid="591" eventid="16" swimtime="00:02:20.36" lane="1" heatid="16002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:08.09" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="592" eventid="32" swimtime="00:01:02.23" lane="5" heatid="32002" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="161" birthdate="2011-01-01" gender="F" lastname="Behrmann" firstname="Fine Erna" license="0">
              <RESULTS>
                <RESULT resultid="593" eventid="1" status="DNS" swimtime="00:00:00.00" lane="2" heatid="1003" />
                <RESULT resultid="594" eventid="15" swimtime="00:02:23.69" lane="7" heatid="15003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:07.38" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="595" eventid="31" status="DNS" swimtime="00:00:00.00" lane="5" heatid="31003" />
                <RESULT resultid="596" eventid="33" status="DNS" swimtime="00:00:00.00" lane="1" heatid="33002" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="162" birthdate="2009-01-01" gender="F" lastname="Henkel" firstname="Friederike" license="0">
              <RESULTS>
                <RESULT resultid="597" eventid="1" swimtime="00:00:26.99" lane="8" heatid="1006" />
                <RESULT resultid="598" eventid="15" swimtime="00:02:19.46" lane="7" heatid="15004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:05.87" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="599" eventid="31" swimtime="00:00:59.23" lane="7" heatid="31004" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="163" birthdate="2008-01-01" gender="M" lastname="Hannemann" firstname="Fynn" license="0">
              <RESULTS>
                <RESULT resultid="600" eventid="14" status="DSQ" swimtime="00:00:58.77" lane="6" heatid="14002" comment="DTG an der Wand bei 50 Meter." />
                <RESULT resultid="601" eventid="16" swimtime="00:01:56.43" lane="8" heatid="16005">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:55.77" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="602" eventid="32" swimtime="00:00:49.83" lane="1" heatid="32007" />
                <RESULT resultid="603" eventid="38" swimtime="00:00:21.28" lane="2" heatid="38004" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="164" birthdate="2009-01-01" gender="M" lastname="Artschwager" firstname="Gustaf" license="0">
              <RESULTS>
                <RESULT resultid="604" eventid="2" swimtime="00:00:25.89" lane="5" heatid="2002" />
                <RESULT resultid="605" eventid="16" swimtime="00:02:07.69" lane="7" heatid="16003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:00.77" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="606" eventid="18" swimtime="00:10:01.57" lane="1" heatid="18002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:05.00" />
                    <SPLIT distance="200" swimtime="00:02:20.47" />
                    <SPLIT distance="300" swimtime="00:03:37.44" />
                    <SPLIT distance="400" swimtime="00:04:54.51" />
                    <SPLIT distance="500" swimtime="00:06:12.39" />
                    <SPLIT distance="600" swimtime="00:07:31.92" />
                    <SPLIT distance="700" swimtime="00:08:50.06" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="607" eventid="32" swimtime="00:00:56.96" lane="4" heatid="32003" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="165" birthdate="1970-01-01" gender="M" lastname="Timpel" firstname="Heiko" license="0">
              <RESULTS>
                <RESULT resultid="608" eventid="2" swimtime="00:00:23.72" lane="8" heatid="2007" />
                <RESULT resultid="609" eventid="14" swimtime="00:00:48.45" lane="8" heatid="14004" />
                <RESULT resultid="610" eventid="20" swimtime="00:04:03.58" lane="4" heatid="20002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:48.30" />
                    <SPLIT distance="200" swimtime="00:01:50.34" />
                    <SPLIT distance="300" swimtime="00:02:56.03" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="611" eventid="32" swimtime="00:00:51.91" lane="8" heatid="32008" />
                <RESULT resultid="612" eventid="38" swimtime="00:00:20.86" lane="2" heatid="38005" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="166" birthdate="2010-01-01" gender="M" lastname="Leipold" firstname="Jakob" license="0">
              <RESULTS>
                <RESULT resultid="613" eventid="2" swimtime="00:00:24.22" lane="7" heatid="2006" />
                <RESULT resultid="614" eventid="14" swimtime="00:00:52.80" lane="5" heatid="14002" />
                <RESULT resultid="615" eventid="16" swimtime="00:01:58.76" lane="6" heatid="16004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:57.28" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="616" eventid="20" swimtime="00:04:55.54" lane="3" heatid="20001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:07.28" />
                    <SPLIT distance="200" swimtime="00:02:23.20" />
                    <SPLIT distance="300" swimtime="00:03:40.59" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="617" eventid="32" swimtime="00:00:53.93" lane="3" heatid="32005" />
                <RESULT resultid="618" eventid="34" swimtime="00:04:26.33" lane="6" heatid="34004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:01.68" />
                    <SPLIT distance="200" swimtime="00:02:11.44" />
                    <SPLIT distance="300" swimtime="00:03:20.72" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="619" eventid="36" swimtime="00:00:23.38" lane="4" heatid="36001" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="167" birthdate="2010-01-01" gender="M" lastname="Hochstein" firstname="Jean Paul" license="0">
              <RESULTS>
                <RESULT resultid="620" eventid="2" swimtime="00:00:24.91" lane="4" heatid="2003" />
                <RESULT resultid="621" eventid="16" swimtime="00:02:13.19" lane="6" heatid="16002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:04.81" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="622" eventid="32" swimtime="00:00:57.03" lane="5" heatid="32003" />
                <RESULT resultid="623" eventid="34" swimtime="00:04:38.96" lane="4" heatid="34002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:05.88" />
                    <SPLIT distance="200" swimtime="00:02:17.92" />
                    <SPLIT distance="300" swimtime="00:03:30.35" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="168" birthdate="2006-01-01" gender="F" lastname="Heinitz" firstname="Leonor" license="0">
              <RESULTS>
                <RESULT resultid="625" eventid="13" swimtime="00:00:50.27" lane="8" heatid="13005" />
                <RESULT resultid="626" eventid="15" swimtime="00:01:58.24" lane="3" heatid="15006">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:56.23" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="627" eventid="31" swimtime="00:00:51.99" lane="3" heatid="31009" />
                <RESULT resultid="628" eventid="33" swimtime="00:04:15.97" lane="3" heatid="33004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:00.47" />
                    <SPLIT distance="200" swimtime="00:02:05.72" />
                    <SPLIT distance="300" swimtime="00:03:12.63" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="629" eventid="37" swimtime="00:00:21.68" lane="2" heatid="37003" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="169" birthdate="2010-01-01" gender="M" lastname="Hochstein" firstname="Maddox Lee" license="0">
              <RESULTS>
                <RESULT resultid="630" eventid="2" swimtime="00:00:27.06" lane="7" heatid="2003" />
                <RESULT resultid="631" eventid="16" swimtime="00:02:17.76" lane="7" heatid="16002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:06.77" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="632" eventid="32" swimtime="00:01:00.21" lane="3" heatid="32002" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="170" birthdate="2006-01-01" gender="M" lastname="Leipold" firstname="Marek" license="0">
              <RESULTS>
                <RESULT resultid="633" eventid="2" swimtime="00:00:16.35" lane="4" heatid="2009" />
                <RESULT resultid="1414" eventid="8" swimtime="00:00:16.54" lane="3" heatid="8001" />
                <RESULT resultid="634" eventid="14" swimtime="00:00:35.28" lane="5" heatid="14006" />
                <RESULT resultid="635" eventid="16" swimtime="00:01:28.53" lane="5" heatid="16008">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:42.99" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1505" eventid="22" swimtime="00:00:35.33" lane="5" heatid="22001" />
                <RESULT resultid="1528" eventid="24" swimtime="00:01:28.67" lane="5" heatid="24001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:42.55" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="636" eventid="32" swimtime="00:00:36.94" lane="4" heatid="32010" />
                <RESULT resultid="637" eventid="38" swimtime="00:00:15.36" lane="5" heatid="38009" />
                <RESULT resultid="1544" eventid="42" swimtime="00:00:37.15" lane="5" heatid="42001" />
                <RESULT resultid="1562" eventid="46" swimtime="00:00:15.42" lane="6" heatid="46001" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="171" birthdate="2009-01-01" gender="F" lastname="Blumenstein" firstname="Martha" license="0">
              <RESULTS>
                <RESULT resultid="638" eventid="1" swimtime="00:00:23.94" lane="7" heatid="1009" />
                <RESULT resultid="639" eventid="3" swimtime="00:18:19.27" lane="5" heatid="3001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:04.07" />
                    <SPLIT distance="200" swimtime="00:02:15.79" />
                    <SPLIT distance="300" swimtime="00:03:28.69" />
                    <SPLIT distance="400" swimtime="00:04:42.45" />
                    <SPLIT distance="500" swimtime="00:05:57.06" />
                    <SPLIT distance="600" swimtime="00:07:11.82" />
                    <SPLIT distance="700" swimtime="00:08:26.44" />
                    <SPLIT distance="800" swimtime="00:09:41.34" />
                    <SPLIT distance="900" swimtime="00:10:55.94" />
                    <SPLIT distance="1000" swimtime="00:12:10.46" />
                    <SPLIT distance="1100" swimtime="00:13:25.07" />
                    <SPLIT distance="1200" swimtime="00:14:39.35" />
                    <SPLIT distance="1300" swimtime="00:15:55.30" />
                    <SPLIT distance="1400" swimtime="00:17:09.25" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="640" eventid="15" swimtime="00:02:06.16" lane="7" heatid="15006">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:01.53" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="641" eventid="17" swimtime="00:09:20.30" lane="1" heatid="17003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:04.44" />
                    <SPLIT distance="200" swimtime="00:02:16.40" />
                    <SPLIT distance="300" swimtime="00:03:29.15" />
                    <SPLIT distance="400" swimtime="00:04:41.38" />
                    <SPLIT distance="500" swimtime="00:05:53.53" />
                    <SPLIT distance="600" swimtime="00:07:05.23" />
                    <SPLIT distance="700" swimtime="00:08:15.69" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="642" eventid="31" swimtime="00:00:53.04" lane="8" heatid="31009" />
                <RESULT resultid="643" eventid="33" swimtime="00:04:32.13" lane="1" heatid="33004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:02.01" />
                    <SPLIT distance="200" swimtime="00:02:13.12" />
                    <SPLIT distance="300" swimtime="00:03:25.90" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="172" birthdate="1978-01-01" gender="M" lastname="Hannemann" firstname="Ronny" license="0">
              <RESULTS>
                <RESULT resultid="644" eventid="14" swimtime="00:00:59.43" lane="8" heatid="14002" />
                <RESULT resultid="645" eventid="32" swimtime="00:00:56.84" lane="4" heatid="32004" />
                <RESULT resultid="646" eventid="38" swimtime="00:00:24.20" lane="8" heatid="38003" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="173" birthdate="1979-01-01" gender="F" lastname="Leipold" firstname="Steffi" license="0">
              <RESULTS>
                <RESULT resultid="647" eventid="1" swimtime="00:00:25.15" lane="4" heatid="1005" />
                <RESULT resultid="648" eventid="15" swimtime="00:02:06.02" lane="7" heatid="15005">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:00.14" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="649" eventid="17" swimtime="00:10:05.00" lane="8" heatid="17003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:04.04" />
                    <SPLIT distance="200" swimtime="00:02:19.71" />
                    <SPLIT distance="300" swimtime="00:03:37.23" />
                    <SPLIT distance="400" swimtime="00:04:53.88" />
                    <SPLIT distance="500" swimtime="00:06:12.54" />
                    <SPLIT distance="600" swimtime="00:07:31.92" />
                    <SPLIT distance="700" swimtime="00:08:50.53" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="650" eventid="31" swimtime="00:00:55.54" lane="2" heatid="31008" />
                <RESULT resultid="651" eventid="33" swimtime="00:04:28.01" lane="7" heatid="33003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:01.19" />
                    <SPLIT distance="200" swimtime="00:02:12.42" />
                    <SPLIT distance="300" swimtime="00:03:22.75" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="652" eventid="37" swimtime="00:00:24.68" lane="6" heatid="37001" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="174" birthdate="1982-01-01" gender="F" lastname="Zitzmann" firstname="Ulrike" license="0">
              <RESULTS>
                <RESULT resultid="653" eventid="1" swimtime="00:00:27.99" lane="7" heatid="1003" />
                <RESULT resultid="655" eventid="5" swimtime="00:01:02.68" lane="3" heatid="5002" />
                <RESULT resultid="656" eventid="39" swimtime="00:00:27.84" lane="1" heatid="39003" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="175" birthdate="1963-01-01" gender="F" lastname="Tiszold" firstname="Ursula" license="0">
              <RESULTS>
                <RESULT resultid="657" eventid="1" swimtime="00:00:31.25" lane="4" heatid="1001" />
                <RESULT resultid="662" eventid="5" swimtime="00:01:10.59" lane="7" heatid="5002" />
                <RESULT resultid="658" eventid="15" swimtime="00:02:39.34" lane="2" heatid="15002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:12.24" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="659" eventid="31" swimtime="00:01:09.11" lane="4" heatid="31002" />
                <RESULT resultid="660" eventid="33" swimtime="00:05:39.91" lane="3" heatid="33001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:16.45" />
                    <SPLIT distance="200" swimtime="00:02:43.29" />
                    <SPLIT distance="300" swimtime="00:04:12.60" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="661" eventid="37" swimtime="00:00:37.54" lane="7" heatid="37001" />
                <RESULT resultid="663" eventid="39" status="DSQ" swimtime="00:00:37.58" lane="4" heatid="39001" comment="Falscher Start." />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY number="1" gender="F" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="562" eventid="11" swimtime="00:08:15.45" lane="4" heatid="11001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:56.30" />
                    <SPLIT distance="200" swimtime="00:01:58.74" />
                    <SPLIT distance="300" swimtime="00:02:58.32" />
                    <SPLIT distance="400" swimtime="00:04:03.25" />
                    <SPLIT distance="500" swimtime="00:05:07.22" />
                    <SPLIT distance="600" swimtime="00:06:20.12" />
                    <SPLIT distance="700" swimtime="00:07:14.98" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="159" number="1" />
                    <RELAYPOSITION athleteid="171" number="2" />
                    <RELAYPOSITION athleteid="162" number="3" />
                    <RELAYPOSITION athleteid="156" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT resultid="563" eventid="48" swimtime="00:03:37.04" lane="8" heatid="48002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:51.41" />
                    <SPLIT distance="200" swimtime="00:01:47.95" />
                    <SPLIT distance="300" swimtime="00:02:46.73" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="156" number="1" />
                    <RELAYPOSITION athleteid="171" number="2" />
                    <RELAYPOSITION athleteid="162" number="3" />
                    <RELAYPOSITION athleteid="159" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" gender="M" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="564" eventid="12" swimtime="00:08:47.22" lane="5" heatid="12001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:04.80" />
                    <SPLIT distance="200" swimtime="00:02:17.76" />
                    <SPLIT distance="300" swimtime="00:03:18.95" />
                    <SPLIT distance="400" swimtime="00:04:27.68" />
                    <SPLIT distance="500" swimtime="00:05:31.81" />
                    <SPLIT distance="600" swimtime="00:06:44.38" />
                    <SPLIT distance="700" swimtime="00:07:43.60" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="160" number="1" />
                    <RELAYPOSITION athleteid="167" number="2" />
                    <RELAYPOSITION athleteid="169" number="3" />
                    <RELAYPOSITION athleteid="166" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT resultid="565" eventid="49" swimtime="00:03:56.66" lane="5" heatid="49001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:58.32" />
                    <SPLIT distance="200" swimtime="00:01:53.95" />
                    <SPLIT distance="300" swimtime="00:02:55.96" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="166" number="1" />
                    <RELAYPOSITION athleteid="167" number="2" />
                    <RELAYPOSITION athleteid="169" number="3" />
                    <RELAYPOSITION athleteid="160" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" gender="X" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="566" eventid="30" swimtime="00:01:39.34" lane="6" heatid="30002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:52.44" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="166" number="1" />
                    <RELAYPOSITION athleteid="161" number="2" />
                    <RELAYPOSITION athleteid="167" number="3" />
                    <RELAYPOSITION athleteid="156" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="2" gender="X" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="567" eventid="47" swimtime="00:03:46.17" lane="3" heatid="47001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:50.53" />
                    <SPLIT distance="200" swimtime="00:01:46.85" />
                    <SPLIT distance="300" swimtime="00:02:50.91" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="165" number="1" />
                    <RELAYPOSITION athleteid="173" number="2" />
                    <RELAYPOSITION athleteid="174" number="3" />
                    <RELAYPOSITION athleteid="172" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="2" gender="X" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="568" eventid="30" swimtime="00:01:33.97" lane="5" heatid="30002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:47.04" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="163" number="1" />
                    <RELAYPOSITION athleteid="171" number="2" />
                    <RELAYPOSITION athleteid="164" number="3" />
                    <RELAYPOSITION athleteid="159" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="4" gender="X" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="1384" eventid="29" status="DSQ" swimtime="00:01:43.24" lane="3" heatid="29001" comment="1. Schwimmer 15m nach dem Start übertaucht.">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:52.44" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="165" number="1" />
                    <RELAYPOSITION athleteid="174" number="2" />
                    <RELAYPOSITION athleteid="172" number="3" />
                    <RELAYPOSITION athleteid="173" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB name="Tauchsportfreunde Dachau e.V." nation="GER" region="34" code="0">
          <ATHLETES>
            <ATHLETE athleteid="208" birthdate="1969-01-01" gender="M" lastname="Sengpiel" firstname="Alexander" license="0">
              <RESULTS>
                <RESULT resultid="801" eventid="18" swimtime="00:10:04.91" lane="3" heatid="18001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:07.40" />
                    <SPLIT distance="200" swimtime="00:02:24.43" />
                    <SPLIT distance="300" swimtime="00:03:42.04" />
                    <SPLIT distance="400" swimtime="00:04:58.89" />
                    <SPLIT distance="500" swimtime="00:06:16.77" />
                    <SPLIT distance="600" swimtime="00:07:35.80" />
                    <SPLIT distance="700" swimtime="00:08:54.25" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="802" eventid="34" swimtime="00:04:47.14" lane="5" heatid="34001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:05.57" />
                    <SPLIT distance="200" swimtime="00:02:21.35" />
                    <SPLIT distance="300" swimtime="00:03:38.01" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="803" eventid="38" swimtime="00:00:22.47" lane="5" heatid="38002" />
                <RESULT resultid="805" eventid="40" swimtime="00:00:26.09" lane="7" heatid="40002" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="TC Chemie Greiz e.V." nation="GER" region="35" code="174117">
          <ATHLETES>
            <ATHLETE athleteid="131" birthdate="2006-01-01" gender="F" lastname="Frauenfelder" firstname="Anneliese" license="0">
              <RESULTS>
                <RESULT resultid="484" eventid="13" swimtime="00:00:48.21" lane="6" heatid="13005" />
                <RESULT resultid="485" eventid="19" swimtime="00:04:12.13" lane="6" heatid="19002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:55.70" />
                    <SPLIT distance="200" swimtime="00:02:00.05" />
                    <SPLIT distance="300" swimtime="00:03:08.64" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="486" eventid="31" swimtime="00:00:48.98" lane="3" heatid="31013" />
                <RESULT resultid="487" eventid="37" swimtime="00:00:21.03" lane="1" heatid="37006" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="132" birthdate="2009-01-01" gender="F" lastname="Naupold" firstname="Celina" license="0">
              <RESULTS>
                <RESULT resultid="488" eventid="1" swimtime="00:00:25.55" lane="6" heatid="1006" />
                <RESULT resultid="489" eventid="13" swimtime="00:00:52.97" lane="6" heatid="13003" />
                <RESULT resultid="490" eventid="31" swimtime="00:00:55.73" lane="3" heatid="31008" />
                <RESULT resultid="491" eventid="37" swimtime="00:00:23.10" lane="7" heatid="37003" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="133" birthdate="2011-01-01" gender="F" lastname="Brendel" firstname="Emma" license="0">
              <RESULTS>
                <RESULT resultid="492" eventid="1" swimtime="00:00:24.78" lane="5" heatid="1004" />
                <RESULT resultid="497" eventid="5" swimtime="00:01:04.22" lane="8" heatid="5003" />
                <RESULT resultid="493" eventid="13" swimtime="00:00:57.71" lane="4" heatid="13002" />
                <RESULT resultid="494" eventid="19" status="DSQ" swimtime="00:05:42.62" lane="1" heatid="19001" comment="Falsche Wende bei 300 Meter.">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:12.73" />
                    <SPLIT distance="200" swimtime="00:02:35.15" />
                    <SPLIT distance="300" swimtime="00:04:04.19" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="495" eventid="31" swimtime="00:00:56.62" lane="2" heatid="31006" />
                <RESULT resultid="496" eventid="35" swimtime="00:00:24.39" lane="6" heatid="35002" />
                <RESULT resultid="1377" eventid="39" swimtime="00:00:29.50" lane="7" heatid="39002" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="134" birthdate="2008-01-01" gender="M" lastname="Lose" firstname="Fabian" license="0">
              <RESULTS>
                <RESULT resultid="498" eventid="2" swimtime="00:00:26.23" lane="3" heatid="2003" />
                <RESULT resultid="500" eventid="6" swimtime="00:00:59.80" lane="4" heatid="6002" />
                <RESULT resultid="499" eventid="34" status="DNS" swimtime="00:00:00.00" lane="2" heatid="34003" />
                <RESULT resultid="501" eventid="40" swimtime="00:00:25.87" lane="2" heatid="40002" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="139" birthdate="2008-01-01" gender="M" lastname="Robenz" firstname="Jean Robin" license="0">
              <RESULTS>
                <RESULT resultid="506" eventid="2" swimtime="00:00:22.48" lane="5" heatid="2005" />
                <RESULT resultid="512" eventid="6" swimtime="00:00:56.05" lane="4" heatid="6001" />
                <RESULT resultid="507" eventid="14" swimtime="00:00:49.47" lane="6" heatid="14001" />
                <RESULT resultid="508" eventid="16" swimtime="00:02:00.13" lane="5" heatid="16003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:57.68" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="510" eventid="34" swimtime="00:04:38.43" lane="7" heatid="34003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:00.97" />
                    <SPLIT distance="200" swimtime="00:02:13.93" />
                    <SPLIT distance="300" swimtime="00:03:30.13" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="511" eventid="38" swimtime="00:00:22.14" lane="5" heatid="38003" />
                <RESULT resultid="513" eventid="40" swimtime="00:00:25.94" lane="1" heatid="40001" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="140" birthdate="2011-01-01" gender="M" lastname="Wyczisk" firstname="Johann" license="0">
              <RESULTS>
                <RESULT resultid="514" eventid="32" swimtime="00:01:06.66" lane="8" heatid="32002" />
                <RESULT resultid="515" eventid="34" swimtime="00:05:07.26" lane="3" heatid="34001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:12.60" />
                    <SPLIT distance="200" swimtime="00:02:30.93" />
                    <SPLIT distance="300" swimtime="00:03:50.94" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="516" eventid="40" swimtime="00:00:33.83" lane="7" heatid="40001" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="141" birthdate="2006-01-01" gender="F" lastname="Löffler" firstname="Johanna" license="0">
              <RESULTS>
                <RESULT resultid="517" eventid="1" swimtime="00:00:23.16" lane="7" heatid="1010" />
                <RESULT resultid="1378" eventid="5" swimtime="00:01:00.37" lane="8" heatid="5004" />
                <RESULT resultid="518" eventid="15" swimtime="00:02:03.12" lane="4" heatid="15007">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:57.14" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="519" eventid="31" swimtime="00:00:54.71" lane="2" heatid="31011" />
                <RESULT resultid="520" eventid="37" swimtime="00:00:20.18" lane="2" heatid="37005" />
                <RESULT resultid="521" eventid="39" swimtime="00:00:27.70" lane="2" heatid="39003" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="142" birthdate="2009-01-01" gender="M" lastname="Heydel" firstname="Linus" license="0">
              <RESULTS>
                <RESULT resultid="522" eventid="2" swimtime="00:00:23.00" lane="3" heatid="2004" />
                <RESULT resultid="523" eventid="14" swimtime="00:00:52.55" lane="7" heatid="14002" />
                <RESULT resultid="524" eventid="20" swimtime="00:04:24.61" lane="4" heatid="20001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:59.89" />
                    <SPLIT distance="200" swimtime="00:02:10.36" />
                    <SPLIT distance="300" swimtime="00:03:21.07" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="525" eventid="34" swimtime="00:04:14.62" lane="8" heatid="34004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:57.71" />
                    <SPLIT distance="200" swimtime="00:02:02.39" />
                    <SPLIT distance="300" swimtime="00:03:10.27" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="526" eventid="38" swimtime="00:00:21.07" lane="8" heatid="38004" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="143" birthdate="2008-01-01" gender="M" lastname="Berger" firstname="Louis" license="0">
              <RESULTS>
                <RESULT resultid="527" eventid="2" swimtime="00:00:19.29" lane="7" heatid="2011" />
                <RESULT resultid="528" eventid="16" swimtime="00:01:42.15" lane="7" heatid="16008">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:47.31" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="529" eventid="32" swimtime="00:00:43.90" lane="1" heatid="32012" />
                <RESULT resultid="530" eventid="38" swimtime="00:00:17.71" lane="8" heatid="38006" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="144" birthdate="2008-01-01" gender="F" lastname="Zschegner" firstname="Lucy" license="0">
              <RESULTS>
                <RESULT resultid="531" eventid="13" swimtime="00:00:52.68" lane="2" heatid="13003" />
                <RESULT resultid="532" eventid="19" swimtime="00:04:25.51" lane="3" heatid="19001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:59.31" />
                    <SPLIT distance="200" swimtime="00:02:09.52" />
                    <SPLIT distance="300" swimtime="00:03:20.47" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="533" eventid="31" swimtime="00:00:56.57" lane="4" heatid="31005" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="145" birthdate="2005-01-01" gender="F" lastname="Kupka" firstname="Miriam" license="0">
              <RESULTS>
                <RESULT resultid="534" eventid="1" swimtime="00:00:20.83" lane="7" heatid="1013" />
                <RESULT resultid="535" eventid="15" swimtime="00:01:45.62" lane="1" heatid="15011">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:50.75" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="536" eventid="31" swimtime="00:00:47.05" lane="1" heatid="31015" />
                <RESULT resultid="537" eventid="33" swimtime="00:03:48.80" lane="2" heatid="33007">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:53.79" />
                    <SPLIT distance="200" swimtime="00:01:51.83" />
                    <SPLIT distance="300" swimtime="00:02:51.92" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="538" eventid="37" swimtime="00:00:19.61" lane="7" heatid="37008" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="146" birthdate="1974-01-01" gender="M" lastname="Kühn" firstname="Ronald" license="0">
              <RESULTS>
                <RESULT resultid="539" eventid="2" swimtime="00:00:24.19" lane="7" heatid="2005" />
                <RESULT resultid="543" eventid="6" swimtime="00:00:57.46" lane="2" heatid="6001" />
                <RESULT resultid="540" eventid="16" swimtime="00:02:03.96" lane="7" heatid="16004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:58.33" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="541" eventid="32" swimtime="00:00:54.54" lane="3" heatid="32006" />
                <RESULT resultid="542" eventid="38" swimtime="00:00:21.64" lane="7" heatid="38004" />
                <RESULT resultid="544" eventid="40" swimtime="00:00:27.01" lane="5" heatid="40001" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="147" birthdate="2011-01-01" gender="F" lastname="Leonhardt" firstname="Ronja" license="0">
              <RESULTS>
                <RESULT resultid="545" eventid="3" swimtime="00:21:34.63" lane="7" heatid="3001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:12.89" />
                    <SPLIT distance="200" swimtime="00:02:38.22" />
                    <SPLIT distance="300" swimtime="00:04:04.95" />
                    <SPLIT distance="400" swimtime="00:05:31.93" />
                    <SPLIT distance="500" swimtime="00:07:00.08" />
                    <SPLIT distance="600" swimtime="00:08:28.45" />
                    <SPLIT distance="700" swimtime="00:09:58.32" />
                    <SPLIT distance="800" swimtime="00:11:28.05" />
                    <SPLIT distance="900" swimtime="00:12:56.65" />
                    <SPLIT distance="1000" swimtime="00:14:24.11" />
                    <SPLIT distance="1100" swimtime="00:15:54.44" />
                    <SPLIT distance="1200" swimtime="00:17:22.90" />
                    <SPLIT distance="1300" swimtime="00:18:51.37" />
                    <SPLIT distance="1400" swimtime="00:20:15.24" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="546" eventid="15" swimtime="00:02:28.57" lane="8" heatid="15002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:11.00" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="547" eventid="17" swimtime="00:10:55.52" lane="5" heatid="17001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:14.86" />
                    <SPLIT distance="200" swimtime="00:02:39.19" />
                    <SPLIT distance="300" swimtime="00:04:04.09" />
                    <SPLIT distance="400" swimtime="00:05:28.33" />
                    <SPLIT distance="500" swimtime="00:06:51.92" />
                    <SPLIT distance="600" swimtime="00:08:16.18" />
                    <SPLIT distance="700" swimtime="00:09:38.77" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="548" eventid="33" swimtime="00:05:20.39" lane="5" heatid="33001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:13.82" />
                    <SPLIT distance="200" swimtime="00:02:37.40" />
                    <SPLIT distance="300" swimtime="00:04:01.97" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="549" eventid="39" swimtime="00:00:31.72" lane="7" heatid="39001" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="148" birthdate="2011-01-01" gender="F" lastname="Klar" firstname="Sophia" license="0">
              <RESULTS>
                <RESULT resultid="550" eventid="1" swimtime="00:00:30.12" lane="2" heatid="1001" />
                <RESULT resultid="554" eventid="5" swimtime="00:01:20.42" lane="3" heatid="5001" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="149" birthdate="2000-01-01" gender="M" lastname="Kupka" firstname="Titus" license="0">
              <RESULTS>
                <RESULT resultid="556" eventid="2" swimtime="00:00:18.61" lane="2" heatid="2011" />
                <RESULT resultid="560" eventid="6" swimtime="00:00:47.08" lane="3" heatid="6004" />
                <RESULT resultid="1419" eventid="8" swimtime="00:00:19.17" lane="8" heatid="8001" />
                <RESULT resultid="557" eventid="14" swimtime="00:00:41.29" lane="3" heatid="14005" />
                <RESULT resultid="558" eventid="32" swimtime="00:00:43.00" lane="7" heatid="32012" />
                <RESULT resultid="559" eventid="38" swimtime="00:00:16.57" lane="6" heatid="38008" />
                <RESULT resultid="561" eventid="40" swimtime="00:00:21.05" lane="4" heatid="40004" />
                <RESULT resultid="1565" eventid="46" swimtime="00:00:16.54" lane="1" heatid="46001" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY number="1" gender="F" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="502" eventid="11" swimtime="00:08:09.74" lane="5" heatid="11002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:53.95" />
                    <SPLIT distance="200" swimtime="00:01:49.02" />
                    <SPLIT distance="300" swimtime="00:02:49.33" />
                    <SPLIT distance="400" swimtime="00:03:58.08" />
                    <SPLIT distance="500" swimtime="00:04:57.83" />
                    <SPLIT distance="600" swimtime="00:06:05.73" />
                    <SPLIT distance="700" swimtime="00:07:03.51" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="145" number="1" />
                    <RELAYPOSITION athleteid="144" number="2" />
                    <RELAYPOSITION athleteid="132" number="3" />
                    <RELAYPOSITION athleteid="141" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" gender="X" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="503" eventid="30" swimtime="00:01:29.96" lane="4" heatid="30002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:47.34" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="144" number="1" />
                    <RELAYPOSITION athleteid="132" number="2" />
                    <RELAYPOSITION athleteid="142" number="3" />
                    <RELAYPOSITION athleteid="143" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" gender="F" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="" />
            <RELAY number="1" gender="F" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="505" eventid="48" swimtime="00:03:22.26" lane="5" heatid="48002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:46.51" />
                    <SPLIT distance="200" swimtime="00:01:38.27" />
                    <SPLIT distance="300" swimtime="00:02:33.23" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="145" number="1" />
                    <RELAYPOSITION athleteid="141" number="2" />
                    <RELAYPOSITION athleteid="144" number="3" />
                    <RELAYPOSITION athleteid="131" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB name="TC Delitzsch" nation="GER" region="20" code="0">
          <ATHLETES>
            <ATHLETE athleteid="194" birthdate="2011-01-01" gender="F" lastname="Schönherr" firstname="Nina" license="0">
              <RESULTS>
                <RESULT resultid="725" eventid="1" swimtime="00:00:25.27" lane="6" heatid="1004" />
                <RESULT resultid="726" eventid="13" swimtime="00:00:56.71" lane="2" heatid="13002" />
                <RESULT resultid="727" eventid="15" swimtime="00:02:11.27" lane="2" heatid="15003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:00.17" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="728" eventid="31" swimtime="00:00:56.69" lane="5" heatid="31007" />
                <RESULT resultid="729" eventid="35" swimtime="00:00:24.65" lane="5" heatid="35001" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="195" birthdate="2011-01-01" gender="M" lastname="Becker" firstname="Pepe Milan" license="0">
              <RESULTS>
                <RESULT resultid="730" eventid="2" swimtime="00:00:26.15" lane="2" heatid="2003" />
                <RESULT resultid="731" eventid="14" swimtime="00:01:05.51" lane="8" heatid="14001" />
                <RESULT resultid="732" eventid="16" swimtime="00:02:14.84" lane="2" heatid="16002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:05.37" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="733" eventid="32" swimtime="00:00:59.90" lane="8" heatid="32003" />
                <RESULT resultid="734" eventid="36" swimtime="00:00:29.95" lane="2" heatid="36001" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="TC fez Berlin" nation="GER" region="21" code="34113000">
          <ATHLETES>
            <ATHLETE athleteid="300" birthdate="2006-01-01" gender="M" lastname="Schlohbohm" firstname="Enrico" license="3411">
              <RESULTS>
                <RESULT resultid="1117" eventid="2" swimtime="00:00:19.24" lane="1" heatid="2011" />
                <RESULT resultid="1118" eventid="14" swimtime="00:00:45.35" lane="1" heatid="14004" />
                <RESULT resultid="1119" eventid="16" swimtime="00:01:45.67" lane="1" heatid="16007">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:49.97" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1120" eventid="32" swimtime="00:00:43.32" lane="7" heatid="32011" />
                <RESULT resultid="1121" eventid="38" status="DNS" swimtime="00:00:00.00" lane="2" heatid="38007" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="301" birthdate="1996-01-01" gender="M" lastname="Schustek" firstname="Fabian" license="0">
              <RESULTS>
                <RESULT resultid="1122" eventid="14" swimtime="00:00:41.73" lane="7" heatid="14004" />
                <RESULT resultid="1123" eventid="16" swimtime="00:01:36.01" lane="2" heatid="16008">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:44.84" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1124" eventid="32" swimtime="00:00:41.06" lane="6" heatid="32010" />
                <RESULT resultid="1125" eventid="38" swimtime="00:00:17.37" lane="1" heatid="38007" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="302" birthdate="2005-01-01" gender="F" lastname="Tesch" firstname="Florentine" license="0">
              <RESULTS>
                <RESULT resultid="1126" eventid="1" swimtime="00:00:19.99" lane="2" heatid="1014" />
                <RESULT resultid="1411" eventid="7" swimtime="00:00:19.63" lane="1" heatid="7001" />
                <RESULT resultid="1127" eventid="9" swimtime="00:16:18.62" lane="3" heatid="9001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:51.16" />
                    <SPLIT distance="200" swimtime="00:01:49.86" />
                    <SPLIT distance="300" swimtime="00:02:51.70" />
                    <SPLIT distance="400" swimtime="00:03:54.79" />
                    <SPLIT distance="500" swimtime="00:04:58.31" />
                    <SPLIT distance="600" swimtime="00:06:03.50" />
                    <SPLIT distance="700" swimtime="00:07:10.23" />
                    <SPLIT distance="800" swimtime="00:08:16.52" />
                    <SPLIT distance="900" swimtime="00:09:23.88" />
                    <SPLIT distance="1000" swimtime="00:10:32.72" />
                    <SPLIT distance="1100" swimtime="00:11:41.93" />
                    <SPLIT distance="1200" swimtime="00:12:49.93" />
                    <SPLIT distance="1300" swimtime="00:13:59.39" />
                    <SPLIT distance="1400" swimtime="00:15:09.74" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1128" eventid="15" swimtime="00:01:48.42" lane="1" heatid="15012">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:50.12" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1129" eventid="25" swimtime="00:07:50.71" lane="1" heatid="25001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:52.06" />
                    <SPLIT distance="200" swimtime="00:01:50.78" />
                    <SPLIT distance="300" swimtime="00:02:51.25" />
                    <SPLIT distance="400" swimtime="00:03:52.48" />
                    <SPLIT distance="500" swimtime="00:04:54.12" />
                    <SPLIT distance="600" swimtime="00:05:54.76" />
                    <SPLIT distance="700" swimtime="00:06:55.30" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1130" eventid="31" swimtime="00:00:46.99" lane="2" heatid="31015" />
                <RESULT resultid="1131" eventid="33" swimtime="00:03:50.74" lane="7" heatid="33007">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:50.70" />
                    <SPLIT distance="200" swimtime="00:01:48.41" />
                    <SPLIT distance="300" swimtime="00:02:49.34" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1386" eventid="37" swimtime="00:00:18.34" lane="3" heatid="37006" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="303" birthdate="2002-01-01" gender="F" lastname="Schikora" firstname="Johanna" license="0">
              <RESULTS>
                <RESULT resultid="1132" eventid="9" swimtime="00:13:29.43" lane="4" heatid="9001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:50.54" />
                    <SPLIT distance="200" swimtime="00:01:41.44" />
                    <SPLIT distance="300" swimtime="00:02:34.07" />
                    <SPLIT distance="400" swimtime="00:03:27.67" />
                    <SPLIT distance="500" swimtime="00:04:21.46" />
                    <SPLIT distance="600" swimtime="00:05:16.14" />
                    <SPLIT distance="700" swimtime="00:06:10.88" />
                    <SPLIT distance="800" swimtime="00:07:05.72" />
                    <SPLIT distance="900" swimtime="00:08:00.60" />
                    <SPLIT distance="1000" swimtime="00:08:55.58" />
                    <SPLIT distance="1100" swimtime="00:09:50.56" />
                    <SPLIT distance="1200" swimtime="00:10:46.15" />
                    <SPLIT distance="1300" swimtime="00:11:40.74" />
                    <SPLIT distance="1400" swimtime="00:12:35.58" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1133" eventid="15" swimtime="00:01:34.13" lane="4" heatid="15011">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:45.98" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1514" eventid="23" swimtime="00:01:32.86" lane="4" heatid="23001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:45.57" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1134" eventid="25" swimtime="00:07:09.34" lane="4" heatid="25001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:51.07" />
                    <SPLIT distance="200" swimtime="00:01:45.38" />
                    <SPLIT distance="300" swimtime="00:02:39.82" />
                    <SPLIT distance="400" swimtime="00:03:34.20" />
                    <SPLIT distance="500" swimtime="00:04:28.88" />
                    <SPLIT distance="600" swimtime="00:05:23.26" />
                    <SPLIT distance="700" swimtime="00:06:17.30" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1135" eventid="31" swimtime="00:00:43.64" lane="5" heatid="31016" />
                <RESULT resultid="1539" eventid="41" swimtime="00:00:43.33" lane="2" heatid="41001" />
                <RESULT resultid="1136" eventid="43" swimtime="00:03:23.88" lane="4" heatid="43001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:48.97" />
                    <SPLIT distance="200" swimtime="00:01:40.48" />
                    <SPLIT distance="300" swimtime="00:02:33.26" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="304" birthdate="2006-01-01" gender="F" lastname="Zobel" firstname="Juliane" license="341100319">
              <RESULTS>
                <RESULT resultid="1137" eventid="1" swimtime="00:00:21.50" lane="7" heatid="1012" />
                <RESULT resultid="1138" eventid="3" swimtime="00:16:40.03" lane="6" heatid="3002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:01.30" />
                    <SPLIT distance="200" swimtime="00:02:08.76" />
                    <SPLIT distance="300" swimtime="00:03:17.51" />
                    <SPLIT distance="400" swimtime="00:04:25.33" />
                    <SPLIT distance="500" swimtime="00:05:34.35" />
                    <SPLIT distance="600" swimtime="00:06:43.87" />
                    <SPLIT distance="700" swimtime="00:07:51.70" />
                    <SPLIT distance="800" swimtime="00:08:59.80" />
                    <SPLIT distance="900" swimtime="00:10:08.22" />
                    <SPLIT distance="1000" swimtime="00:11:16.15" />
                    <SPLIT distance="1100" swimtime="00:12:23.59" />
                    <SPLIT distance="1200" swimtime="00:13:31.12" />
                    <SPLIT distance="1300" swimtime="00:14:37.32" />
                    <SPLIT distance="1400" swimtime="00:15:41.60" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1139" eventid="15" swimtime="00:01:48.22" lane="5" heatid="15009">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:52.22" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1140" eventid="17" swimtime="00:08:21.88" lane="3" heatid="17004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:57.64" />
                    <SPLIT distance="200" swimtime="00:02:01.58" />
                    <SPLIT distance="300" swimtime="00:03:06.63" />
                    <SPLIT distance="400" swimtime="00:04:11.73" />
                    <SPLIT distance="500" swimtime="00:05:16.65" />
                    <SPLIT distance="600" swimtime="00:06:21.23" />
                    <SPLIT distance="700" swimtime="00:07:24.47" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1141" eventid="31" swimtime="00:00:47.79" lane="5" heatid="31013" />
                <RESULT resultid="1142" eventid="37" swimtime="00:00:20.15" lane="4" heatid="37003" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="305" birthdate="2005-01-01" gender="F" lastname="Gawenda" firstname="Lara" license="0">
              <RESULTS>
                <RESULT resultid="1143" eventid="1" swimtime="00:00:18.85" lane="4" heatid="1013" />
                <RESULT resultid="1404" eventid="7" swimtime="00:00:18.97" lane="4" heatid="7001" />
                <RESULT resultid="1144" eventid="15" swimtime="00:01:36.37" lane="5" heatid="15011">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:46.58" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1516" eventid="23" swimtime="00:01:36.40" lane="3" heatid="23001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:46.25" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1145" eventid="31" swimtime="00:00:42.78" lane="4" heatid="31015" />
                <RESULT resultid="1146" eventid="37" swimtime="00:00:18.02" lane="4" heatid="37006" />
                <RESULT resultid="1536" eventid="41" swimtime="00:00:46.21" lane="5" heatid="41001" />
                <RESULT resultid="1555" eventid="45" swimtime="00:00:18.03" lane="2" heatid="45001" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="306" birthdate="2007-01-01" gender="F" lastname="Schikora" firstname="Luise" license="0">
              <RESULTS>
                <RESULT resultid="1147" eventid="1" swimtime="00:00:21.94" lane="1" heatid="1012" />
                <RESULT resultid="1148" eventid="15" swimtime="00:01:50.80" lane="7" heatid="15008">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:52.41" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1149" eventid="31" swimtime="00:00:46.88" lane="4" heatid="31012" />
                <RESULT resultid="1150" eventid="37" swimtime="00:00:19.19" lane="7" heatid="37004" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="307" birthdate="2007-01-01" gender="F" lastname="Rüdiger" firstname="Marielena" license="0">
              <RESULTS>
                <RESULT resultid="1151" eventid="1" swimtime="00:00:26.65" lane="5" heatid="1006" />
                <RESULT resultid="1152" eventid="15" swimtime="00:02:06.48" lane="5" heatid="15005">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:01.98" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1153" eventid="31" swimtime="00:00:57.98" lane="4" heatid="31007" />
                <RESULT resultid="1154" eventid="33" swimtime="00:04:46.19" lane="8" heatid="33003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:08.78" />
                    <SPLIT distance="200" swimtime="00:02:25.47" />
                    <SPLIT distance="300" swimtime="00:03:39.53" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1155" eventid="37" swimtime="00:00:23.28" lane="5" heatid="37001" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="308" birthdate="2000-01-01" gender="F" lastname="Teichler" firstname="Maxi" license="0">
              <RESULTS>
                <RESULT resultid="1156" eventid="13" swimtime="00:00:53.50" lane="8" heatid="13006" />
                <RESULT resultid="1157" eventid="31" swimtime="00:00:53.82" lane="8" heatid="31011" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="309" birthdate="2008-01-01" gender="F" lastname="Sunagatova" firstname="Milana" license="0">
              <RESULTS>
                <RESULT resultid="1158" eventid="1" swimtime="00:00:20.85" lane="2" heatid="1013" />
                <RESULT resultid="1159" eventid="15" swimtime="00:01:43.67" lane="7" heatid="15010">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:49.99" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1160" eventid="25" swimtime="00:08:08.86" lane="7" heatid="25001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:54.01" />
                    <SPLIT distance="200" swimtime="00:01:55.55" />
                    <SPLIT distance="300" swimtime="00:02:58.52" />
                    <SPLIT distance="400" swimtime="00:04:01.21" />
                    <SPLIT distance="500" swimtime="00:05:04.15" />
                    <SPLIT distance="600" swimtime="00:06:07.36" />
                    <SPLIT distance="700" swimtime="00:07:10.37" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1161" eventid="31" swimtime="00:00:46.23" lane="7" heatid="31017" />
                <RESULT resultid="1162" eventid="43" swimtime="00:03:51.01" lane="7" heatid="43001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:53.03" />
                    <SPLIT distance="200" swimtime="00:01:52.21" />
                    <SPLIT distance="300" swimtime="00:02:52.82" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="310" birthdate="2006-01-01" gender="F" lastname="Ahnert" firstname="Paula" license="0">
              <RESULTS>
                <RESULT resultid="1163" eventid="1" swimtime="00:00:20.77" lane="6" heatid="1010" />
                <RESULT resultid="1164" eventid="3" swimtime="00:15:41.03" lane="4" heatid="3001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:53.69" />
                    <SPLIT distance="200" swimtime="00:01:52.88" />
                    <SPLIT distance="300" swimtime="00:02:54.94" />
                    <SPLIT distance="400" swimtime="00:03:57.99" />
                    <SPLIT distance="500" swimtime="00:05:01.47" />
                    <SPLIT distance="600" swimtime="00:06:05.70" />
                    <SPLIT distance="700" swimtime="00:07:09.87" />
                    <SPLIT distance="800" swimtime="00:08:13.82" />
                    <SPLIT distance="900" swimtime="00:09:17.76" />
                    <SPLIT distance="1000" swimtime="00:10:21.99" />
                    <SPLIT distance="1100" swimtime="00:11:25.86" />
                    <SPLIT distance="1200" swimtime="00:12:30.38" />
                    <SPLIT distance="1300" swimtime="00:13:34.92" />
                    <SPLIT distance="1400" swimtime="00:14:38.98" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1165" eventid="15" swimtime="00:01:43.16" lane="8" heatid="15009">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:49.07" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1166" eventid="17" swimtime="00:08:16.64" lane="8" heatid="17005">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:53.57" />
                    <SPLIT distance="200" swimtime="00:01:52.90" />
                    <SPLIT distance="300" swimtime="00:02:54.90" />
                    <SPLIT distance="400" swimtime="00:03:58.21" />
                    <SPLIT distance="500" swimtime="00:05:03.63" />
                    <SPLIT distance="600" swimtime="00:06:08.83" />
                    <SPLIT distance="700" swimtime="00:07:13.12" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1167" eventid="31" swimtime="00:00:43.58" lane="4" heatid="31008" />
                <RESULT resultid="1168" eventid="33" status="DNS" swimtime="00:00:00.00" lane="3" heatid="33005" />
                <RESULT resultid="1538" eventid="41" swimtime="00:00:44.11" lane="6" heatid="41001" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="311" birthdate="1996-01-01" gender="M" lastname="Wegner" firstname="Pit" license="0">
              <RESULTS>
                <RESULT resultid="1169" eventid="38" swimtime="00:00:20.28" lane="4" heatid="38005" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="312" birthdate="2002-01-01" gender="M" lastname="Lebeau" firstname="Remy" license="0">
              <RESULTS>
                <RESULT resultid="1170" eventid="2" swimtime="00:00:19.24" lane="6" heatid="2010" />
                <RESULT resultid="1385" eventid="14" swimtime="00:00:38.23" lane="6" heatid="14005" />
                <RESULT resultid="1503" eventid="22" status="WDR" swimtime="00:00:00.00" lane="0" heatid="22000" />
                <RESULT resultid="1172" eventid="28" swimtime="00:03:00.68" lane="7" heatid="28001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:41.70" />
                    <SPLIT distance="200" swimtime="00:01:27.62" />
                    <SPLIT distance="300" swimtime="00:02:15.24" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1173" eventid="32" swimtime="00:00:42.20" lane="5" heatid="32010" />
                <RESULT resultid="1174" eventid="44" swimtime="00:03:17.61" lane="5" heatid="44001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:45.98" />
                    <SPLIT distance="200" swimtime="00:01:35.92" />
                    <SPLIT distance="300" swimtime="00:02:26.90" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="313" birthdate="2006-01-01" gender="M" lastname="Patge" firstname="Rufus" license="3411">
              <RESULTS>
                <RESULT resultid="1175" eventid="10" swimtime="00:16:41.62" lane="2" heatid="10001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:58.22" />
                    <SPLIT distance="200" swimtime="00:02:01.33" />
                    <SPLIT distance="300" swimtime="00:03:09.77" />
                    <SPLIT distance="400" swimtime="00:04:14.09" />
                    <SPLIT distance="500" swimtime="00:05:18.96" />
                    <SPLIT distance="600" swimtime="00:06:26.23" />
                    <SPLIT distance="700" swimtime="00:07:32.73" />
                    <SPLIT distance="800" swimtime="00:08:40.49" />
                    <SPLIT distance="900" swimtime="00:09:48.86" />
                    <SPLIT distance="1000" swimtime="00:10:59.92" />
                    <SPLIT distance="1100" swimtime="00:12:09.69" />
                    <SPLIT distance="1200" swimtime="00:13:18.17" />
                    <SPLIT distance="1300" swimtime="00:14:27.60" />
                    <SPLIT distance="1400" swimtime="00:15:34.40" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1176" eventid="16" swimtime="00:01:45.58" lane="7" heatid="16007">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:50.36" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1177" eventid="26" swimtime="00:08:02.99" lane="1" heatid="26001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:53.16" />
                    <SPLIT distance="200" swimtime="00:01:53.42" />
                    <SPLIT distance="300" swimtime="00:02:56.33" />
                    <SPLIT distance="400" swimtime="00:03:59.18" />
                    <SPLIT distance="500" swimtime="00:05:01.33" />
                    <SPLIT distance="600" swimtime="00:06:03.16" />
                    <SPLIT distance="700" swimtime="00:07:03.60" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1178" eventid="28" swimtime="00:03:46.61" lane="1" heatid="28001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:52.38" />
                    <SPLIT distance="200" swimtime="00:01:49.63" />
                    <SPLIT distance="300" swimtime="00:02:48.59" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1179" eventid="34" swimtime="00:03:48.41" lane="3" heatid="34006">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:51.47" />
                    <SPLIT distance="200" swimtime="00:01:50.61" />
                    <SPLIT distance="300" swimtime="00:02:50.18" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="314" birthdate="2005-01-01" gender="F" lastname="Hoffmann" firstname="Zoe" license="0">
              <RESULTS>
                <RESULT resultid="1180" eventid="1" swimtime="00:00:23.93" lane="6" heatid="1008" />
                <RESULT resultid="1181" eventid="31" swimtime="00:00:55.05" lane="7" heatid="31009" />
                <RESULT resultid="1182" eventid="37" swimtime="00:00:22.74" lane="1" heatid="37003" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="375" birthdate="1995-01-01" gender="M" lastname="Willruth" firstname="Tim" license="0" />
          </ATHLETES>
          <RELAYS>
            <RELAY number="1" gender="M" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="1109" eventid="12" swimtime="00:06:47.13" lane="3" heatid="12002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:47.25" />
                    <SPLIT distance="200" swimtime="00:01:43.78" />
                    <SPLIT distance="300" swimtime="00:02:32.68" />
                    <SPLIT distance="400" swimtime="00:03:28.85" />
                    <SPLIT distance="500" swimtime="00:04:17.29" />
                    <SPLIT distance="600" swimtime="00:05:11.85" />
                    <SPLIT distance="700" swimtime="00:05:55.75" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="300" number="1" />
                    <RELAYPOSITION athleteid="313" number="2" />
                    <RELAYPOSITION athleteid="375" number="3" />
                    <RELAYPOSITION athleteid="301" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT resultid="1110" eventid="49" swimtime="00:02:50.78" lane="5" heatid="49002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:42.40" />
                    <SPLIT distance="200" swimtime="00:01:26.28" />
                    <SPLIT distance="300" swimtime="00:02:10.95" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="300" number="1" />
                    <RELAYPOSITION athleteid="375" number="2" />
                    <RELAYPOSITION athleteid="313" number="3" />
                    <RELAYPOSITION athleteid="301" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" gender="F" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="1111" eventid="11" swimtime="00:06:36.41" lane="4" heatid="11003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:46.99" />
                    <SPLIT distance="200" swimtime="00:01:37.65" />
                    <SPLIT distance="300" swimtime="00:02:22.87" />
                    <SPLIT distance="400" swimtime="00:03:10.95" />
                    <SPLIT distance="500" swimtime="00:03:58.10" />
                    <SPLIT distance="600" swimtime="00:04:53.30" />
                    <SPLIT distance="700" swimtime="00:05:40.72" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="305" number="1" />
                    <RELAYPOSITION athleteid="303" number="2" />
                    <RELAYPOSITION athleteid="310" number="3" />
                    <RELAYPOSITION athleteid="302" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT resultid="1112" eventid="48" swimtime="00:02:53.22" lane="4" heatid="48003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:43.13" />
                    <SPLIT distance="200" swimtime="00:01:26.12" />
                    <SPLIT distance="300" swimtime="00:02:09.03" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="305" number="1" />
                    <RELAYPOSITION athleteid="303" number="2" />
                    <RELAYPOSITION athleteid="310" number="3" />
                    <RELAYPOSITION athleteid="302" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" gender="X" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="1113" eventid="30" swimtime="00:01:15.59" lane="8" heatid="30004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:38.63" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="305" number="1" />
                    <RELAYPOSITION athleteid="303" number="2" />
                    <RELAYPOSITION athleteid="301" number="3" />
                    <RELAYPOSITION athleteid="375" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="2" gender="F" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="1114" eventid="11" swimtime="00:07:40.17" lane="1" heatid="11003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:50.52" />
                    <SPLIT distance="200" swimtime="00:01:46.79" />
                    <SPLIT distance="300" swimtime="00:02:36.83" />
                    <SPLIT distance="400" swimtime="00:03:38.06" />
                    <SPLIT distance="500" swimtime="00:04:42.22" />
                    <SPLIT distance="600" swimtime="00:05:46.56" />
                    <SPLIT distance="700" swimtime="00:06:39.80" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="309" number="1" />
                    <RELAYPOSITION athleteid="306" number="2" />
                    <RELAYPOSITION athleteid="307" number="3" />
                    <RELAYPOSITION athleteid="304" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT resultid="1115" eventid="48" swimtime="00:03:17.99" lane="4" heatid="48002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:48.15" />
                    <SPLIT distance="200" swimtime="00:01:35.90" />
                    <SPLIT distance="300" swimtime="00:02:31.26" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="304" number="1" />
                    <RELAYPOSITION athleteid="306" number="2" />
                    <RELAYPOSITION athleteid="307" number="3" />
                    <RELAYPOSITION athleteid="309" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="2" gender="X" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="1116" eventid="30" swimtime="00:01:20.13" lane="6" heatid="30003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:38.67" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="310" number="1" />
                    <RELAYPOSITION athleteid="300" number="2" />
                    <RELAYPOSITION athleteid="313" number="3" />
                    <RELAYPOSITION athleteid="304" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB name="TC Marzahn e.V." nation="GER" region="21" code="0">
          <ATHLETES>
            <ATHLETE athleteid="216" birthdate="2010-01-01" gender="F" lastname="Liedloff" firstname="Amelie" license="0">
              <RESULTS>
                <RESULT resultid="821" eventid="1" swimtime="00:00:22.98" lane="4" heatid="1011" />
                <RESULT resultid="822" eventid="3" swimtime="00:19:17.35" lane="3" heatid="3001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:04.51" />
                    <SPLIT distance="200" swimtime="00:02:18.03" />
                    <SPLIT distance="300" swimtime="00:03:39.52" />
                    <SPLIT distance="400" swimtime="00:04:59.52" />
                    <SPLIT distance="500" swimtime="00:06:22.44" />
                    <SPLIT distance="600" swimtime="00:07:43.25" />
                    <SPLIT distance="700" swimtime="00:09:03.99" />
                    <SPLIT distance="800" swimtime="00:10:26.97" />
                    <SPLIT distance="900" swimtime="00:11:49.62" />
                    <SPLIT distance="1000" swimtime="00:13:12.27" />
                    <SPLIT distance="1100" swimtime="00:14:29.52" />
                    <SPLIT distance="1200" swimtime="00:15:51.01" />
                    <SPLIT distance="1300" swimtime="00:17:02.97" />
                    <SPLIT distance="1400" swimtime="00:18:10.83" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="823" eventid="15" swimtime="00:01:58.16" lane="5" heatid="15007">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:54.03" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="824" eventid="17" swimtime="00:09:50.90" lane="8" heatid="17004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:07.38" />
                    <SPLIT distance="200" swimtime="00:02:22.99" />
                    <SPLIT distance="300" swimtime="00:03:40.11" />
                    <SPLIT distance="400" swimtime="00:04:57.09" />
                    <SPLIT distance="500" swimtime="00:06:15.45" />
                    <SPLIT distance="600" swimtime="00:07:34.30" />
                    <SPLIT distance="700" swimtime="00:08:45.52" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="825" eventid="31" swimtime="00:00:52.59" lane="4" heatid="31011" />
                <RESULT resultid="826" eventid="33" swimtime="00:04:24.40" lane="1" heatid="33006">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:00.56" />
                    <SPLIT distance="200" swimtime="00:02:09.69" />
                    <SPLIT distance="300" swimtime="00:03:19.52" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="217" birthdate="1965-01-01" gender="M" lastname="Ritzer" firstname="Andre" license="0">
              <RESULTS>
                <RESULT resultid="827" eventid="2" swimtime="00:00:27.39" lane="8" heatid="2004" />
                <RESULT resultid="831" eventid="6" swimtime="00:01:01.74" lane="5" heatid="6002" />
                <RESULT resultid="828" eventid="16" swimtime="00:02:14.16" lane="5" heatid="16002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:01.59" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="829" eventid="32" swimtime="00:01:00.25" lane="1" heatid="32004" />
                <RESULT resultid="830" eventid="38" swimtime="00:00:23.98" lane="1" heatid="38003" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="218" birthdate="2010-01-01" gender="F" lastname="Kempe" firstname="Anna" license="0">
              <RESULTS>
                <RESULT resultid="832" eventid="1" swimtime="00:00:26.97" lane="1" heatid="1003" />
                <RESULT resultid="833" eventid="15" swimtime="00:02:23.46" lane="8" heatid="15003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:12.80" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="834" eventid="31" swimtime="00:01:01.70" lane="2" heatid="31005" />
                <RESULT resultid="835" eventid="39" swimtime="00:00:31.24" lane="3" heatid="39001" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="219" birthdate="1977-01-01" gender="F" lastname="Lopez" firstname="Annett" license="0">
              <RESULTS>
                <RESULT resultid="836" eventid="1" swimtime="00:00:25.51" lane="1" heatid="1007" />
                <RESULT resultid="837" eventid="15" swimtime="00:02:02.18" lane="2" heatid="15006">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:58.34" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="838" eventid="17" swimtime="00:09:41.41" lane="2" heatid="17003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:04.59" />
                    <SPLIT distance="200" swimtime="00:02:16.40" />
                    <SPLIT distance="300" swimtime="00:03:29.31" />
                    <SPLIT distance="400" swimtime="00:04:43.38" />
                    <SPLIT distance="500" swimtime="00:05:57.83" />
                    <SPLIT distance="600" swimtime="00:07:13.96" />
                    <SPLIT distance="700" swimtime="00:08:29.98" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="839" eventid="31" swimtime="00:00:56.60" lane="7" heatid="31008" />
                <RESULT resultid="840" eventid="33" swimtime="00:04:31.79" lane="4" heatid="33003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:01.26" />
                    <SPLIT distance="200" swimtime="00:02:10.76" />
                    <SPLIT distance="300" swimtime="00:03:22.04" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="220" birthdate="2008-01-01" gender="F" lastname="Demmrich" firstname="Ella" license="0">
              <RESULTS>
                <RESULT resultid="841" eventid="1" swimtime="00:00:27.86" lane="4" heatid="1004" />
                <RESULT resultid="847" eventid="5" swimtime="00:01:01.21" lane="6" heatid="5003" />
                <RESULT resultid="842" eventid="15" swimtime="00:02:04.66" lane="3" heatid="15005">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:59.30" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="843" eventid="17" swimtime="00:09:42.10" lane="3" heatid="17002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:02.76" />
                    <SPLIT distance="200" swimtime="00:02:14.90" />
                    <SPLIT distance="300" swimtime="00:03:30.04" />
                    <SPLIT distance="400" swimtime="00:04:45.75" />
                    <SPLIT distance="500" swimtime="00:06:01.86" />
                    <SPLIT distance="600" swimtime="00:07:17.60" />
                    <SPLIT distance="700" swimtime="00:08:31.58" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="844" eventid="31" swimtime="00:00:58.52" lane="6" heatid="31006" />
                <RESULT resultid="845" eventid="33" swimtime="00:04:38.10" lane="6" heatid="33002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:03.36" />
                    <SPLIT distance="200" swimtime="00:02:15.51" />
                    <SPLIT distance="300" swimtime="00:03:29.35" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="846" eventid="37" swimtime="00:00:24.93" lane="2" heatid="37001" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="221" birthdate="2009-01-01" gender="M" lastname="Kupke" firstname="Emil" license="0">
              <RESULTS>
                <RESULT resultid="848" eventid="2" swimtime="00:00:24.94" lane="6" heatid="2004" />
                <RESULT resultid="849" eventid="16" swimtime="00:02:09.63" lane="3" heatid="16002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:02.25" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="850" eventid="32" swimtime="00:00:56.09" lane="7" heatid="32004" />
                <RESULT resultid="851" eventid="34" swimtime="00:04:53.41" lane="6" heatid="34002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:07.84" />
                    <SPLIT distance="200" swimtime="00:02:22.97" />
                    <SPLIT distance="300" swimtime="00:03:40.48" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="852" eventid="38" swimtime="00:00:23.64" lane="2" heatid="38002" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="222" birthdate="2004-01-01" gender="F" lastname="May" firstname="Emilie" license="0">
              <RESULTS>
                <RESULT resultid="853" eventid="1" swimtime="00:00:22.27" lane="1" heatid="1011" />
                <RESULT resultid="855" eventid="5" swimtime="00:00:54.64" lane="5" heatid="5004" />
                <RESULT resultid="1381" eventid="31" swimtime="00:00:47.36" lane="5" heatid="31011" />
                <RESULT resultid="854" eventid="37" swimtime="00:00:19.85" lane="5" heatid="37004" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="223" birthdate="2009-01-01" gender="M" lastname="Müller" firstname="Erik" license="0">
              <RESULTS>
                <RESULT resultid="856" eventid="2" swimtime="00:00:25.94" lane="7" heatid="2002" />
                <RESULT resultid="858" eventid="6" swimtime="00:01:00.35" lane="3" heatid="6001" />
                <RESULT resultid="857" eventid="32" swimtime="00:01:00.18" lane="2" heatid="32002" />
                <RESULT resultid="859" eventid="40" swimtime="00:00:26.47" lane="6" heatid="40001" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="224" birthdate="2005-01-01" gender="M" lastname="Kwauka" firstname="Kevin" license="0">
              <RESULTS>
                <RESULT resultid="860" eventid="2" swimtime="00:00:19.52" lane="1" heatid="2010" />
                <RESULT resultid="861" eventid="14" swimtime="00:00:45.81" lane="8" heatid="14006" />
                <RESULT resultid="862" eventid="32" swimtime="00:00:46.57" lane="4" heatid="32008" />
                <RESULT resultid="863" eventid="38" swimtime="00:00:18.33" lane="8" heatid="38008" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="225" birthdate="2005-01-01" gender="F" lastname="Eweleit" firstname="Laura" license="0">
              <RESULTS>
                <RESULT resultid="864" eventid="1" swimtime="00:00:20.76" lane="3" heatid="1013" />
                <RESULT resultid="865" eventid="9" status="DSQ" swimtime="00:14:47.67" lane="7" heatid="9001" comment="Tauchzüge außerhalb der 15m Zone.">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:54.68" />
                    <SPLIT distance="200" swimtime="00:01:52.70" />
                    <SPLIT distance="300" swimtime="00:02:51.63" />
                    <SPLIT distance="400" swimtime="00:03:51.28" />
                    <SPLIT distance="500" swimtime="00:04:51.03" />
                    <SPLIT distance="600" swimtime="00:05:51.19" />
                    <SPLIT distance="700" swimtime="00:06:51.31" />
                    <SPLIT distance="800" swimtime="00:07:50.22" />
                    <SPLIT distance="900" swimtime="00:08:50.29" />
                    <SPLIT distance="1000" swimtime="00:09:50.56" />
                    <SPLIT distance="1100" swimtime="00:10:50.39" />
                    <SPLIT distance="1200" swimtime="00:11:50.97" />
                    <SPLIT distance="1300" swimtime="00:12:51.06" />
                    <SPLIT distance="1400" swimtime="00:13:50.88" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="866" eventid="15" swimtime="00:01:42.33" lane="3" heatid="15011">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:49.04" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="867" eventid="25" swimtime="00:07:42.15" lane="3" heatid="25001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:53.01" />
                    <SPLIT distance="200" swimtime="00:01:50.88" />
                    <SPLIT distance="300" swimtime="00:02:50.80" />
                    <SPLIT distance="400" swimtime="00:03:49.65" />
                    <SPLIT distance="500" swimtime="00:04:49.35" />
                    <SPLIT distance="600" swimtime="00:05:48.56" />
                    <SPLIT distance="700" swimtime="00:06:46.47" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="868" eventid="31" swimtime="00:00:44.94" lane="2" heatid="31017" />
                <RESULT resultid="870" eventid="37" swimtime="00:00:18.96" lane="6" heatid="37008" />
                <RESULT resultid="1534" eventid="41" status="WDR" swimtime="00:00:00.00" lane="0" heatid="41000" />
                <RESULT resultid="869" eventid="43" swimtime="00:03:38.90" lane="6" heatid="43001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:51.57" />
                    <SPLIT distance="200" swimtime="00:01:46.72" />
                    <SPLIT distance="300" swimtime="00:02:43.78" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="226" birthdate="2010-01-01" gender="F" lastname="Haupt" firstname="Lena" license="0">
              <RESULTS>
                <RESULT resultid="871" eventid="1" swimtime="00:00:23.90" lane="3" heatid="1007" />
                <RESULT resultid="875" eventid="5" swimtime="00:00:57.06" lane="4" heatid="5003" />
                <RESULT resultid="872" eventid="15" swimtime="00:01:58.56" lane="2" heatid="15007">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:55.75" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="873" eventid="17" swimtime="00:09:32.18" lane="5" heatid="17002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:06.45" />
                    <SPLIT distance="200" swimtime="00:02:18.98" />
                    <SPLIT distance="300" swimtime="00:03:32.45" />
                    <SPLIT distance="400" swimtime="00:04:46.20" />
                    <SPLIT distance="500" swimtime="00:05:59.60" />
                    <SPLIT distance="600" swimtime="00:07:12.49" />
                    <SPLIT distance="700" swimtime="00:08:24.46" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="874" eventid="31" swimtime="00:00:55.06" lane="5" heatid="31008" />
                <RESULT resultid="876" eventid="39" swimtime="00:00:26.12" lane="3" heatid="39003" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="227" birthdate="2011-01-01" gender="F" lastname="Eweleit" firstname="Lenja" license="0">
              <RESULTS>
                <RESULT resultid="877" eventid="1" swimtime="00:00:25.83" lane="7" heatid="1005" />
                <RESULT resultid="878" eventid="15" swimtime="00:02:07.92" lane="8" heatid="15005">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:02.69" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="879" eventid="17" swimtime="00:09:39.25" lane="7" heatid="17002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:07.67" />
                    <SPLIT distance="200" swimtime="00:02:20.79" />
                    <SPLIT distance="300" swimtime="00:03:34.54" />
                    <SPLIT distance="400" swimtime="00:04:48.30" />
                    <SPLIT distance="500" swimtime="00:06:02.68" />
                    <SPLIT distance="600" swimtime="00:07:17.39" />
                    <SPLIT distance="700" swimtime="00:08:31.59" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="880" eventid="31" swimtime="00:00:59.42" lane="5" heatid="31006" />
                <RESULT resultid="881" eventid="33" swimtime="00:04:39.66" lane="1" heatid="33003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:06.21" />
                    <SPLIT distance="200" swimtime="00:02:19.26" />
                    <SPLIT distance="300" swimtime="00:03:31.50" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="228" birthdate="2005-01-01" gender="F" lastname="Marleen Reinbach" firstname="Lilly" license="0">
              <RESULTS>
                <RESULT resultid="882" eventid="1" swimtime="00:00:22.81" lane="7" heatid="1011" />
                <RESULT resultid="886" eventid="5" swimtime="00:00:59.66" lane="5" heatid="5003" />
                <RESULT resultid="883" eventid="13" swimtime="00:00:47.67" lane="3" heatid="13004" />
                <RESULT resultid="884" eventid="31" swimtime="00:00:51.46" lane="5" heatid="31012" />
                <RESULT resultid="885" eventid="37" swimtime="00:00:21.33" lane="4" heatid="37004" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="229" birthdate="2001-01-01" gender="M" lastname="Lopez" firstname="Marvin" license="0">
              <RESULTS>
                <RESULT resultid="887" eventid="2" swimtime="00:00:19.45" lane="2" heatid="2010" />
                <RESULT resultid="888" eventid="16" swimtime="00:01:40.04" lane="2" heatid="16006">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:47.16" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="889" eventid="32" status="DSQ" swimtime="00:00:00.00" lane="1" heatid="32011" comment="Aufgegeben nach 60 Meter." />
                <RESULT resultid="890" eventid="38" swimtime="00:00:17.79" lane="7" heatid="38008" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="230" birthdate="1971-01-01" gender="M" lastname="Tech" firstname="Matthias" license="0">
              <RESULTS>
                <RESULT resultid="891" eventid="2" swimtime="00:00:22.98" lane="1" heatid="2007" />
                <RESULT resultid="1379" eventid="6" swimtime="00:00:56.31" lane="6" heatid="6003" />
                <RESULT resultid="892" eventid="32" swimtime="00:00:53.50" lane="2" heatid="32006" />
                <RESULT resultid="893" eventid="38" swimtime="00:00:20.21" lane="7" heatid="38005" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="231" birthdate="1982-01-01" gender="F" lastname="Heilek" firstname="Sarah" license="0">
              <RESULTS>
                <RESULT resultid="894" eventid="31" swimtime="00:01:04.78" lane="6" heatid="31003" />
                <RESULT resultid="895" eventid="39" swimtime="00:00:31.05" lane="6" heatid="39001" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="232" birthdate="2007-01-01" gender="F" lastname="Götz" firstname="Zoe" license="0">
              <RESULTS>
                <RESULT resultid="896" eventid="1" swimtime="00:00:22.24" lane="3" heatid="1011" />
                <RESULT resultid="903" eventid="5" swimtime="00:00:57.92" lane="6" heatid="5004" />
                <RESULT resultid="897" eventid="13" swimtime="00:00:47.73" lane="1" heatid="13007" />
                <RESULT resultid="898" eventid="15" swimtime="00:01:57.86" lane="4" heatid="15008">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:58.17" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="899" eventid="19" swimtime="00:04:38.39" lane="7" heatid="19001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:03.63" />
                    <SPLIT distance="200" swimtime="00:02:14.37" />
                    <SPLIT distance="300" swimtime="00:03:28.24" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="900" eventid="31" swimtime="00:00:48.91" lane="1" heatid="31013" />
                <RESULT resultid="901" eventid="33" swimtime="00:04:18.95" lane="8" heatid="33006">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:59.32" />
                    <SPLIT distance="200" swimtime="00:02:05.67" />
                    <SPLIT distance="300" swimtime="00:03:14.32" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="902" eventid="37" swimtime="00:00:20.33" lane="3" heatid="37004" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY number="2" gender="M" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="812" eventid="12" status="DNS" swimtime="00:00:00.00" lane="7" heatid="12002">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="229" number="1" />
                    <RELAYPOSITION athleteid="224" number="2" />
                    <RELAYPOSITION athleteid="223" number="3" />
                    <RELAYPOSITION athleteid="221" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT resultid="813" eventid="49" swimtime="00:03:26.22" lane="1" heatid="49002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:42.48" />
                    <SPLIT distance="200" swimtime="00:01:28.80" />
                    <SPLIT distance="300" swimtime="00:02:26.22" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="229" number="1" />
                    <RELAYPOSITION athleteid="224" number="2" />
                    <RELAYPOSITION athleteid="223" number="3" />
                    <RELAYPOSITION athleteid="221" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="3" gender="F" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="814" eventid="11" swimtime="00:08:33.32" lane="3" heatid="11002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:55.97" />
                    <SPLIT distance="200" swimtime="00:02:00.56" />
                    <SPLIT distance="300" swimtime="00:02:57.74" />
                    <SPLIT distance="400" swimtime="00:04:00.51" />
                    <SPLIT distance="500" swimtime="00:05:04.66" />
                    <SPLIT distance="600" swimtime="00:06:09.46" />
                    <SPLIT distance="700" swimtime="00:07:15.89" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="216" number="1" />
                    <RELAYPOSITION athleteid="226" number="2" />
                    <RELAYPOSITION athleteid="227" number="3" />
                    <RELAYPOSITION athleteid="218" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT resultid="816" eventid="48" swimtime="00:03:46.93" lane="2" heatid="48002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:52.47" />
                    <SPLIT distance="200" swimtime="00:01:48.10" />
                    <SPLIT distance="300" swimtime="00:02:46.83" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="216" number="1" />
                    <RELAYPOSITION athleteid="226" number="2" />
                    <RELAYPOSITION athleteid="227" number="3" />
                    <RELAYPOSITION athleteid="218" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" gender="F" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="815" eventid="11" swimtime="00:07:17.80" lane="7" heatid="11003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:49.92" />
                    <SPLIT distance="200" swimtime="00:01:44.17" />
                    <SPLIT distance="300" swimtime="00:02:34.03" />
                    <SPLIT distance="400" swimtime="00:03:30.43" />
                    <SPLIT distance="500" swimtime="00:04:23.53" />
                    <SPLIT distance="600" swimtime="00:05:21.29" />
                    <SPLIT distance="700" swimtime="00:06:16.29" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="225" number="1" />
                    <RELAYPOSITION athleteid="222" number="2" />
                    <RELAYPOSITION athleteid="228" number="3" />
                    <RELAYPOSITION athleteid="232" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT resultid="817" eventid="48" swimtime="00:03:11.09" lane="1" heatid="48003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:44.93" />
                    <SPLIT distance="200" swimtime="00:01:32.01" />
                    <SPLIT distance="300" swimtime="00:02:22.31" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="225" number="1" />
                    <RELAYPOSITION athleteid="222" number="2" />
                    <RELAYPOSITION athleteid="228" number="3" />
                    <RELAYPOSITION athleteid="232" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="4" gender="X" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="818" eventid="30" swimtime="00:01:19.44" lane="2" heatid="30004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:38.45" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="229" number="1" />
                    <RELAYPOSITION athleteid="224" number="2" />
                    <RELAYPOSITION athleteid="222" number="3" />
                    <RELAYPOSITION athleteid="225" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="5" gender="X" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="819" eventid="30" swimtime="00:01:37.57" lane="3" heatid="30002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:48.47" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="226" number="1" />
                    <RELAYPOSITION athleteid="221" number="2" />
                    <RELAYPOSITION athleteid="223" number="3" />
                    <RELAYPOSITION athleteid="216" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="6" gender="X" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="820" eventid="47" swimtime="00:03:52.87" lane="6" heatid="47001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:56.05" />
                    <SPLIT distance="200" swimtime="00:01:48.59" />
                    <SPLIT distance="300" swimtime="00:02:48.74" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="219" number="1" />
                    <RELAYPOSITION athleteid="230" number="2" />
                    <RELAYPOSITION athleteid="217" number="3" />
                    <RELAYPOSITION athleteid="231" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB name="TC Nautilus Mitterteich" nation="GER" region="34" code="24135">
          <ATHLETES>
            <ATHLETE athleteid="9" birthdate="1992-01-01" gender="F" lastname="Schaller" firstname="Christin" license="0">
              <RESULTS>
                <RESULT resultid="46" eventid="1" swimtime="00:00:28.18" lane="8" heatid="1004" />
                <RESULT resultid="47" eventid="13" swimtime="00:00:59.20" lane="5" heatid="13002" />
                <RESULT resultid="1380" eventid="19" swimtime="00:05:13.29" lane="6" heatid="19001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:06.29" />
                    <SPLIT distance="200" swimtime="00:02:27.35" />
                    <SPLIT distance="300" swimtime="00:03:53.42" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="49" eventid="31" swimtime="00:01:02.26" lane="8" heatid="31005" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="TC submarin Pößneck" nation="GER" region="35" code="174116000">
          <ATHLETES>
            <ATHLETE athleteid="275" birthdate="2005-01-01" gender="F" lastname="Heinze" firstname="Charlotte" license="0">
              <RESULTS>
                <RESULT resultid="1046" eventid="13" swimtime="00:00:45.76" lane="3" heatid="13005" />
                <RESULT resultid="1047" eventid="19" swimtime="00:04:01.96" lane="4" heatid="19002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:53.20" />
                    <SPLIT distance="200" swimtime="00:01:53.13" />
                    <SPLIT distance="300" swimtime="00:02:54.67" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1048" eventid="37" swimtime="00:00:19.44" lane="2" heatid="37007" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="276" birthdate="2007-01-01" gender="F" lastname="Näther" firstname="Emilia" license="0">
              <RESULTS>
                <RESULT resultid="1049" eventid="1" swimtime="00:00:20.43" lane="7" heatid="1015" />
                <RESULT resultid="1050" eventid="31" swimtime="00:00:46.35" lane="8" heatid="31014" />
                <RESULT resultid="1051" eventid="37" swimtime="00:00:18.98" lane="1" heatid="37007" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="277" birthdate="2011-01-01" gender="F" lastname="Müller" firstname="Emily" license="0">
              <RESULTS>
                <RESULT resultid="1054" eventid="15" swimtime="00:02:23.26" lane="7" heatid="15002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:08.84" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1055" eventid="17" status="DSQ" swimtime="00:00:00.00" lane="3" heatid="17001" comment="Aufgegeben nach 600 Meter.">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:16.75" />
                    <SPLIT distance="200" swimtime="00:02:41.83" />
                    <SPLIT distance="300" swimtime="00:04:08.56" />
                    <SPLIT distance="400" swimtime="00:05:35.62" />
                    <SPLIT distance="500" swimtime="00:07:00.57" />
                    <SPLIT distance="600" swimtime="00:08:28.33" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1057" eventid="31" swimtime="00:01:03.21" lane="5" heatid="31002" />
                <RESULT resultid="1058" eventid="33" swimtime="00:05:04.16" lane="4" heatid="33001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:10.92" />
                    <SPLIT distance="200" swimtime="00:02:29.08" />
                    <SPLIT distance="300" swimtime="00:03:49.64" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1059" eventid="35" swimtime="00:00:27.70" lane="3" heatid="35001" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="278" birthdate="2005-01-01" gender="F" lastname="Rattke" firstname="Ninette" license="0">
              <RESULTS>
                <RESULT resultid="1060" eventid="3" swimtime="00:18:05.64" lane="2" heatid="3002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:01.36" />
                    <SPLIT distance="200" swimtime="00:02:10.07" />
                    <SPLIT distance="300" swimtime="00:03:20.89" />
                    <SPLIT distance="400" swimtime="00:04:31.82" />
                    <SPLIT distance="500" swimtime="00:05:43.91" />
                    <SPLIT distance="600" swimtime="00:06:57.61" />
                    <SPLIT distance="700" swimtime="00:08:11.93" />
                    <SPLIT distance="800" swimtime="00:09:26.39" />
                    <SPLIT distance="900" swimtime="00:10:42.95" />
                    <SPLIT distance="1000" swimtime="00:11:57.58" />
                    <SPLIT distance="1100" swimtime="00:13:14.73" />
                    <SPLIT distance="1200" swimtime="00:14:32.89" />
                    <SPLIT distance="1300" swimtime="00:15:48.73" />
                    <SPLIT distance="1400" swimtime="00:17:01.49" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1061" eventid="13" swimtime="00:00:47.03" lane="2" heatid="13005" />
                <RESULT resultid="1062" eventid="17" swimtime="00:09:08.51" lane="4" heatid="17004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:58.66" />
                    <SPLIT distance="200" swimtime="00:02:06.78" />
                    <SPLIT distance="300" swimtime="00:03:16.54" />
                    <SPLIT distance="400" swimtime="00:04:28.63" />
                    <SPLIT distance="500" swimtime="00:05:40.80" />
                    <SPLIT distance="600" swimtime="00:06:53.30" />
                    <SPLIT distance="700" swimtime="00:08:04.29" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1063" eventid="19" swimtime="00:04:10.69" lane="2" heatid="19002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:54.49" />
                    <SPLIT distance="200" swimtime="00:01:59.67" />
                    <SPLIT distance="300" swimtime="00:03:07.71" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1064" eventid="31" swimtime="00:00:48.19" lane="3" heatid="31014" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="281" birthdate="2010-01-01" gender="F" lastname="Matthes" firstname="Sophie" license="0">
              <RESULTS>
                <RESULT resultid="1073" eventid="1" swimtime="00:00:25.53" lane="1" heatid="1005" />
                <RESULT resultid="1074" eventid="13" swimtime="00:00:57.46" lane="3" heatid="13001" />
                <RESULT resultid="1075" eventid="15" swimtime="00:02:23.76" lane="1" heatid="15003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:08.66" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1076" eventid="31" swimtime="00:00:57.70" lane="7" heatid="31005" />
                <RESULT resultid="1078" eventid="35" swimtime="00:00:25.28" lane="2" heatid="35002" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="376" birthdate="2011-01-01" gender="M" lastname="Knoblich" firstname="Paul" license="0" />
            <ATHLETE athleteid="377" birthdate="2011-01-01" gender="M" lastname="Rattke" firstname="Carlos" license="0" />
          </ATHLETES>
          <RELAYS>
            <RELAY number="1" gender="X" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="1072" eventid="30" swimtime="00:01:58.11" lane="7" heatid="30002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:05.57" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="376" number="1" />
                    <RELAYPOSITION athleteid="377" number="2" />
                    <RELAYPOSITION athleteid="277" number="3" />
                    <RELAYPOSITION athleteid="281" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB name="The Netherlands" nation="NED" region="0" code="0">
          <ATHLETES>
            <ATHLETE athleteid="64" birthdate="1991-01-01" gender="M" lastname="Cornelissen" firstname="Roelant" license="9259164">
              <RESULTS>
                <RESULT resultid="208" eventid="2" status="DSQ" swimtime="00:00:21.60" lane="6" heatid="2007" comment="Falscher Start." />
                <RESULT resultid="211" eventid="6" swimtime="00:00:52.22" lane="7" heatid="6004" />
                <RESULT resultid="209" eventid="32" swimtime="00:00:50.98" lane="8" heatid="32007" />
                <RESULT resultid="210" eventid="38" swimtime="00:00:18.72" lane="5" heatid="38005" />
                <RESULT resultid="212" eventid="40" swimtime="00:00:22.77" lane="4" heatid="40003" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="65" birthdate="2008-01-01" gender="F" lastname="van der Geest" firstname="Silke" license="9261622">
              <RESULTS>
                <RESULT resultid="213" eventid="1" swimtime="00:00:25.40" lane="7" heatid="1007" />
                <RESULT resultid="216" eventid="5" swimtime="00:01:04.07" lane="4" heatid="5002" />
                <RESULT resultid="214" eventid="15" swimtime="00:02:14.00" lane="4" heatid="15004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:59.80" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="215" eventid="31" swimtime="00:00:57.06" lane="6" heatid="31007" />
                <RESULT resultid="217" eventid="39" swimtime="00:00:28.41" lane="3" heatid="39002" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="66" birthdate="2001-01-01" gender="M" lastname="van Diepen" firstname="Wouter" license="9013676">
              <RESULTS>
                <RESULT resultid="220" eventid="6" swimtime="00:00:49.52" lane="5" heatid="6004" />
                <RESULT resultid="218" eventid="26" swimtime="00:07:25.84" lane="2" heatid="26001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:50.68" />
                    <SPLIT distance="200" swimtime="00:01:46.12" />
                    <SPLIT distance="300" swimtime="00:02:42.86" />
                    <SPLIT distance="400" swimtime="00:03:40.43" />
                    <SPLIT distance="500" swimtime="00:04:37.64" />
                    <SPLIT distance="600" swimtime="00:05:34.61" />
                    <SPLIT distance="700" swimtime="00:06:31.20" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="219" eventid="32" swimtime="00:00:44.09" lane="8" heatid="32012" />
                <RESULT resultid="221" eventid="40" swimtime="00:00:23.16" lane="1" heatid="40004" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="TSC Rostock 1957" nation="GER" region="22" code="0">
          <ATHLETES>
            <ATHLETE athleteid="327" birthdate="2008-01-01" gender="F" lastname="Kellermann" firstname="Alma" license="0">
              <RESULTS>
                <RESULT resultid="1229" eventid="1" swimtime="00:00:19.47" lane="5" heatid="1014" />
                <RESULT resultid="1406" eventid="7" status="DSQ" swimtime="00:00:19.59" lane="3" heatid="7001" comment="Falscher Start." />
                <RESULT resultid="1230" eventid="13" swimtime="00:00:40.64" lane="8" heatid="13001" />
                <RESULT resultid="1231" eventid="15" swimtime="00:01:42.11" lane="7" heatid="15011">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:51.33" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1495" eventid="21" swimtime="00:00:41.80" lane="3" heatid="21001" />
                <RESULT resultid="1520" eventid="23" swimtime="00:01:48.33" lane="1" heatid="23001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:51.39" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1232" eventid="27" swimtime="00:03:34.67" lane="3" heatid="27001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:50.58" />
                    <SPLIT distance="200" swimtime="00:01:45.90" />
                    <SPLIT distance="300" swimtime="00:02:44.02" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1233" eventid="31" swimtime="00:00:44.50" lane="3" heatid="31016" />
                <RESULT resultid="1234" eventid="37" swimtime="00:00:18.15" lane="3" heatid="37008" />
                <RESULT resultid="1542" eventid="41" swimtime="00:00:44.96" lane="8" heatid="41001" />
                <RESULT resultid="1558" eventid="45" swimtime="00:00:18.20" lane="8" heatid="45001" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="328" birthdate="2008-01-01" gender="F" lastname="Schröder" firstname="Alma" license="0">
              <RESULTS>
                <RESULT resultid="1235" eventid="1" swimtime="00:00:27.76" lane="3" heatid="1006" />
                <RESULT resultid="1236" eventid="15" swimtime="00:02:22.66" lane="1" heatid="15005">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:04.36" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1237" eventid="31" status="DNS" swimtime="00:00:00.00" lane="3" heatid="31005" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="329" birthdate="2010-01-01" gender="F" lastname="Timmer" firstname="Anna Fee" license="0">
              <RESULTS>
                <RESULT resultid="1238" eventid="1" swimtime="00:00:30.83" lane="3" heatid="1001" />
                <RESULT resultid="1240" eventid="5" swimtime="00:01:08.52" lane="6" heatid="5002" />
                <RESULT resultid="1239" eventid="31" swimtime="00:01:07.01" lane="4" heatid="31001" />
                <RESULT resultid="1241" eventid="39" swimtime="00:00:29.63" lane="2" heatid="39002" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="330" birthdate="2011-01-01" gender="F" lastname="Meyer" firstname="Anna Lena" license="0">
              <RESULTS>
                <RESULT resultid="1242" eventid="1" swimtime="00:00:31.32" lane="6" heatid="1001" />
                <RESULT resultid="1244" eventid="5" status="DSQ" swimtime="00:01:21.02" lane="4" heatid="5001" comment="Falsche Ausrüstung." />
                <RESULT resultid="1243" eventid="31" swimtime="00:01:09.48" lane="8" heatid="31002" />
                <RESULT resultid="1245" eventid="39" swimtime="00:00:31.66" lane="8" heatid="39002" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="331" birthdate="2011-01-01" gender="M" lastname="Mende" firstname="Bruno" license="0">
              <RESULTS>
                <RESULT resultid="1246" eventid="2" swimtime="00:00:32.59" lane="1" heatid="2001" />
                <RESULT resultid="1247" eventid="32" swimtime="00:01:18.40" lane="6" heatid="32001" />
                <RESULT resultid="1248" eventid="36" swimtime="00:00:32.27" lane="7" heatid="36001" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="332" birthdate="2009-01-01" gender="F" lastname="Mende" firstname="Carla" license="0">
              <RESULTS>
                <RESULT resultid="1249" eventid="1" swimtime="00:00:28.07" lane="6" heatid="1002" />
                <RESULT resultid="1250" eventid="13" status="DSQ" swimtime="00:01:03.67" lane="7" heatid="13001" comment="DTG an der Anschlagmatte bei 100 Meter." />
                <RESULT resultid="1251" eventid="31" swimtime="00:01:04.58" lane="7" heatid="31002" />
                <RESULT resultid="1252" eventid="37" swimtime="00:00:25.38" lane="3" heatid="37001" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="333" birthdate="2006-01-01" gender="F" lastname="Mencke" firstname="Elisa" license="0">
              <RESULTS>
                <RESULT resultid="1253" eventid="3" swimtime="00:17:23.95" lane="5" heatid="3002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:03.55" />
                    <SPLIT distance="200" swimtime="00:02:11.64" />
                    <SPLIT distance="300" swimtime="00:03:20.59" />
                    <SPLIT distance="400" swimtime="00:04:30.10" />
                    <SPLIT distance="500" swimtime="00:05:40.55" />
                    <SPLIT distance="600" swimtime="00:06:50.60" />
                    <SPLIT distance="700" swimtime="00:08:01.13" />
                    <SPLIT distance="800" swimtime="00:09:11.59" />
                    <SPLIT distance="900" swimtime="00:10:21.46" />
                    <SPLIT distance="1000" swimtime="00:11:32.35" />
                    <SPLIT distance="1100" swimtime="00:12:43.11" />
                    <SPLIT distance="1200" swimtime="00:13:54.24" />
                    <SPLIT distance="1300" swimtime="00:15:06.34" />
                    <SPLIT distance="1400" swimtime="00:16:15.99" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1254" eventid="17" swimtime="00:08:26.96" lane="3" heatid="17005">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:59.33" />
                    <SPLIT distance="200" swimtime="00:02:03.36" />
                    <SPLIT distance="300" swimtime="00:03:08.29" />
                    <SPLIT distance="400" swimtime="00:04:13.03" />
                    <SPLIT distance="500" swimtime="00:05:17.36" />
                    <SPLIT distance="600" swimtime="00:06:22.06" />
                    <SPLIT distance="700" swimtime="00:07:25.66" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1255" eventid="31" swimtime="00:00:50.05" lane="2" heatid="31013" />
                <RESULT resultid="1256" eventid="33" swimtime="00:04:03.61" lane="5" heatid="33006">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:57.60" />
                    <SPLIT distance="200" swimtime="00:02:00.36" />
                    <SPLIT distance="300" swimtime="00:03:03.47" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="334" birthdate="2011-01-01" gender="F" lastname="Drews" firstname="Elsa" license="0">
              <RESULTS>
                <RESULT resultid="1257" eventid="15" status="DSQ" swimtime="00:03:34.05" lane="3" heatid="15001" comment="Bei 120m an der Leine festgehalten. Ab 100m Schnorchel nicht zur Atmung benutzt.">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:18.99" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1258" eventid="31" swimtime="00:01:15.85" lane="5" heatid="31001" />
                <RESULT resultid="1259" eventid="39" swimtime="00:00:31.42" lane="1" heatid="39002" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="335" birthdate="2004-01-01" gender="M" lastname="Warning" firstname="Emil" license="0">
              <RESULTS>
                <RESULT resultid="1260" eventid="2" swimtime="00:00:18.71" lane="6" heatid="2009" />
                <RESULT resultid="1261" eventid="14" swimtime="00:00:43.38" lane="2" heatid="14006" />
                <RESULT resultid="1262" eventid="38" swimtime="00:00:17.73" lane="1" heatid="38009" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="336" birthdate="2004-01-01" gender="M" lastname="Malchow" firstname="Finn" license="0">
              <RESULTS>
                <RESULT resultid="1263" eventid="16" swimtime="00:01:29.96" lane="5" heatid="16006">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:43.46" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1529" eventid="24" swimtime="00:01:31.45" lane="3" heatid="24001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:43.70" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1264" eventid="32" swimtime="00:00:40.93" lane="6" heatid="32011" />
                <RESULT resultid="1266" eventid="38" swimtime="00:00:17.53" lane="8" heatid="38005" />
                <RESULT resultid="1550" eventid="42" swimtime="00:00:41.00" lane="8" heatid="42001" />
                <RESULT resultid="1265" eventid="44" swimtime="00:03:25.68" lane="6" heatid="44001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:47.13" />
                    <SPLIT distance="200" swimtime="00:01:39.05" />
                    <SPLIT distance="300" swimtime="00:02:33.00" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="337" birthdate="2008-01-01" gender="F" lastname="Behrend" firstname="Freya" license="0">
              <RESULTS>
                <RESULT resultid="1267" eventid="1" swimtime="00:00:22.70" lane="3" heatid="1009" />
                <RESULT resultid="1268" eventid="13" swimtime="00:00:47.55" lane="1" heatid="13005" />
                <RESULT resultid="1269" eventid="15" swimtime="00:01:58.94" lane="2" heatid="15008">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:57.79" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1270" eventid="31" swimtime="00:00:56.35" lane="8" heatid="31012" />
                <RESULT resultid="1271" eventid="37" swimtime="00:00:21.62" lane="3" heatid="37002" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="338" birthdate="2010-01-01" gender="F" lastname="Buch" firstname="Freya" license="0">
              <RESULTS>
                <RESULT resultid="1272" eventid="1" swimtime="00:00:26.45" lane="5" heatid="1003" />
                <RESULT resultid="1387" eventid="13" swimtime="00:01:01.32" lane="2" heatid="13001" />
                <RESULT resultid="1274" eventid="31" swimtime="00:01:01.10" lane="6" heatid="31005" />
                <RESULT resultid="1275" eventid="33" swimtime="00:04:37.55" lane="2" heatid="33003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:05.78" />
                    <SPLIT distance="200" swimtime="00:02:18.45" />
                    <SPLIT distance="300" swimtime="00:03:31.75" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="339" birthdate="2009-01-01" gender="F" lastname="Kuntz" firstname="Friederike" license="0">
              <RESULTS>
                <RESULT resultid="1276" eventid="1" swimtime="00:00:26.55" lane="4" heatid="1007" />
                <RESULT resultid="1277" eventid="15" swimtime="00:02:12.08" lane="6" heatid="15005">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:05.32" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1278" eventid="33" swimtime="00:04:36.51" lane="8" heatid="33004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:04.50" />
                    <SPLIT distance="200" swimtime="00:02:16.42" />
                    <SPLIT distance="300" swimtime="00:03:27.81" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="340" birthdate="2011-01-01" gender="M" lastname="Behrend" firstname="Gustav" license="0">
              <RESULTS>
                <RESULT resultid="1279" eventid="2" status="DNS" swimtime="00:00:00.00" lane="2" heatid="2001" />
                <RESULT resultid="1280" eventid="16" status="DNS" swimtime="00:00:00.00" lane="6" heatid="16001" />
                <RESULT resultid="1281" eventid="32" status="DNS" swimtime="00:00:00.00" lane="5" heatid="32001" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="341" birthdate="2009-01-01" gender="F" lastname="Gelbricht" firstname="Hedi" license="0">
              <RESULTS>
                <RESULT resultid="1282" eventid="1" swimtime="00:00:24.18" lane="3" heatid="1005" />
                <RESULT resultid="1283" eventid="13" swimtime="00:00:55.26" lane="1" heatid="13003" />
                <RESULT resultid="1284" eventid="15" swimtime="00:02:03.69" lane="1" heatid="15006">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:59.57" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1285" eventid="31" swimtime="00:00:55.65" lane="6" heatid="31008" />
                <RESULT resultid="1286" eventid="33" swimtime="00:04:23.77" lane="2" heatid="33004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:01.60" />
                    <SPLIT distance="200" swimtime="00:02:09.26" />
                    <SPLIT distance="300" swimtime="00:03:18.41" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="342" birthdate="2011-01-01" gender="F" lastname="Beerbaum" firstname="Isabella" license="0">
              <RESULTS>
                <RESULT resultid="1287" eventid="1" swimtime="00:00:30.69" lane="7" heatid="1001" />
                <RESULT resultid="1288" eventid="15" swimtime="00:02:31.87" lane="5" heatid="15001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:09.54" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1289" eventid="31" swimtime="00:01:09.49" lane="1" heatid="31002" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="343" birthdate="2009-01-01" gender="M" lastname="Wippler" firstname="Jannik" license="0">
              <RESULTS>
                <RESULT resultid="1290" eventid="2" swimtime="00:00:28.79" lane="1" heatid="2002" />
                <RESULT resultid="1291" eventid="18" swimtime="00:10:41.52" lane="7" heatid="18002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:09.64" />
                    <SPLIT distance="200" swimtime="00:02:32.01" />
                    <SPLIT distance="300" swimtime="00:03:55.54" />
                    <SPLIT distance="400" swimtime="00:05:18.77" />
                    <SPLIT distance="500" swimtime="00:06:43.06" />
                    <SPLIT distance="600" swimtime="00:08:06.65" />
                    <SPLIT distance="700" swimtime="00:09:29.85" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1292" eventid="34" swimtime="00:05:07.09" lane="2" heatid="34002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:09.68" />
                    <SPLIT distance="200" swimtime="00:02:30.70" />
                    <SPLIT distance="300" swimtime="00:03:52.62" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1293" eventid="38" swimtime="00:00:27.48" lane="5" heatid="38001" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="344" birthdate="2010-01-01" gender="F" lastname="Reichardt" firstname="Jula" license="0">
              <RESULTS>
                <RESULT resultid="1294" eventid="1" swimtime="00:00:27.20" lane="7" heatid="1004" />
                <RESULT resultid="1295" eventid="15" swimtime="00:02:12.92" lane="1" heatid="15004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:03.99" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1296" eventid="17" swimtime="00:10:01.67" lane="4" heatid="17002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:07.80" />
                    <SPLIT distance="200" swimtime="00:02:24.21" />
                    <SPLIT distance="300" swimtime="00:03:41.61" />
                    <SPLIT distance="400" swimtime="00:04:59.06" />
                    <SPLIT distance="500" swimtime="00:06:16.27" />
                    <SPLIT distance="600" swimtime="00:07:35.13" />
                    <SPLIT distance="700" swimtime="00:08:51.50" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1297" eventid="33" swimtime="00:04:50.35" lane="6" heatid="33003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:07.83" />
                    <SPLIT distance="200" swimtime="00:02:23.26" />
                    <SPLIT distance="300" swimtime="00:03:39.86" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="345" birthdate="2011-01-01" gender="M" lastname="Schröder" firstname="Laurent" license="0">
              <RESULTS>
                <RESULT resultid="1298" eventid="2" swimtime="00:00:30.16" lane="3" heatid="2001" />
                <RESULT resultid="1299" eventid="16" swimtime="00:02:37.58" lane="3" heatid="16001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:19.08" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1300" eventid="32" swimtime="00:01:08.69" lane="4" heatid="32001" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="346" birthdate="1998-01-01" gender="F" lastname="Dethloff" firstname="Lisa" license="0">
              <RESULTS>
                <RESULT resultid="1301" eventid="15" swimtime="00:01:42.17" lane="6" heatid="15010">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:49.43" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1521" eventid="23" swimtime="00:01:48.79" lane="8" heatid="23001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:52.17" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1302" eventid="27" swimtime="00:03:25.00" lane="5" heatid="27001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:48.83" />
                    <SPLIT distance="200" swimtime="00:01:40.06" />
                    <SPLIT distance="300" swimtime="00:02:32.37" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="347" birthdate="2010-01-01" gender="M" lastname="Koslov" firstname="Luis" license="0">
              <RESULTS>
                <RESULT resultid="1303" eventid="2" swimtime="00:00:25.81" lane="1" heatid="2003" />
                <RESULT resultid="1304" eventid="14" swimtime="00:00:58.41" lane="2" heatid="14001" />
                <RESULT resultid="1305" eventid="16" swimtime="00:02:10.43" lane="2" heatid="16003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:03.90" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1306" eventid="32" swimtime="00:00:58.22" lane="2" heatid="32004" />
                <RESULT resultid="1307" eventid="34" swimtime="00:04:42.49" lane="6" heatid="34003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:05.93" />
                    <SPLIT distance="200" swimtime="00:02:20.18" />
                    <SPLIT distance="300" swimtime="00:03:34.19" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="348" birthdate="2006-01-01" gender="F" lastname="Stemmler" firstname="Marit" license="0">
              <RESULTS>
                <RESULT resultid="1308" eventid="1" status="DSQ" swimtime="00:00:20.63" lane="5" heatid="1011" comment="Falscher Start." />
                <RESULT resultid="1309" eventid="15" swimtime="00:01:48.80" lane="8" heatid="15010">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:51.44" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1310" eventid="31" swimtime="00:00:47.29" lane="1" heatid="31016" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="349" birthdate="2010-01-01" gender="F" lastname="Peetz" firstname="Marthe" license="0">
              <RESULTS>
                <RESULT resultid="1311" eventid="1" swimtime="00:00:30.16" lane="3" heatid="1002" />
                <RESULT resultid="1313" eventid="5" swimtime="00:01:10.83" lane="2" heatid="5002" />
                <RESULT resultid="1312" eventid="31" swimtime="00:01:11.40" lane="3" heatid="31002" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="350" birthdate="2008-01-01" gender="F" lastname="Drewelow" firstname="Mia" license="0">
              <RESULTS>
                <RESULT resultid="1314" eventid="1" swimtime="00:00:28.43" lane="4" heatid="1002" />
                <RESULT resultid="1315" eventid="15" swimtime="00:02:16.00" lane="5" heatid="15003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:05.93" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1316" eventid="31" swimtime="00:01:03.62" lane="2" heatid="31004" />
                <RESULT resultid="1317" eventid="33" swimtime="00:04:46.32" lane="3" heatid="33002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:07.49" />
                    <SPLIT distance="200" swimtime="00:02:20.92" />
                    <SPLIT distance="300" swimtime="00:03:35.70" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="351" birthdate="2007-01-01" gender="F" lastname="Hecht" firstname="Paula" license="0">
              <RESULTS>
                <RESULT resultid="1318" eventid="1" swimtime="00:00:22.57" lane="5" heatid="1009" />
                <RESULT resultid="1319" eventid="31" swimtime="00:00:50.97" lane="3" heatid="31012" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="352" birthdate="1955-01-01" gender="M" lastname="Szadkowski" firstname="Peter" license="0">
              <RESULTS>
                <RESULT resultid="1320" eventid="18" swimtime="00:11:41.73" lane="6" heatid="18001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:07.37" />
                    <SPLIT distance="200" swimtime="00:02:34.66" />
                    <SPLIT distance="300" swimtime="00:04:04.94" />
                    <SPLIT distance="400" swimtime="00:05:36.69" />
                    <SPLIT distance="500" swimtime="00:07:09.02" />
                    <SPLIT distance="600" swimtime="00:08:40.93" />
                    <SPLIT distance="700" swimtime="00:10:12.10" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1321" eventid="32" swimtime="00:01:04.61" lane="1" heatid="32002" />
                <RESULT resultid="1322" eventid="38" swimtime="00:00:27.49" lane="3" heatid="38001" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="353" birthdate="2009-01-01" gender="M" lastname="Riegmann" firstname="Timo" license="0">
              <RESULTS>
                <RESULT resultid="1323" eventid="10" swimtime="00:17:13.97" lane="7" heatid="10001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:05.72" />
                    <SPLIT distance="200" swimtime="00:02:14.67" />
                    <SPLIT distance="300" swimtime="00:03:25.96" />
                    <SPLIT distance="400" swimtime="00:04:38.73" />
                    <SPLIT distance="500" swimtime="00:05:50.57" />
                    <SPLIT distance="600" swimtime="00:07:02.39" />
                    <SPLIT distance="700" swimtime="00:08:15.14" />
                    <SPLIT distance="800" swimtime="00:09:26.72" />
                    <SPLIT distance="900" swimtime="00:10:36.86" />
                    <SPLIT distance="1000" swimtime="00:11:45.72" />
                    <SPLIT distance="1100" swimtime="00:12:53.58" />
                    <SPLIT distance="1200" swimtime="00:14:01.22" />
                    <SPLIT distance="1300" swimtime="00:15:07.39" />
                    <SPLIT distance="1400" swimtime="00:16:12.37" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1324" eventid="18" swimtime="00:08:56.21" lane="4" heatid="18003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:04.74" />
                    <SPLIT distance="200" swimtime="00:02:13.77" />
                    <SPLIT distance="300" swimtime="00:03:24.30" />
                    <SPLIT distance="400" swimtime="00:04:33.59" />
                    <SPLIT distance="500" swimtime="00:05:42.15" />
                    <SPLIT distance="600" swimtime="00:06:49.61" />
                    <SPLIT distance="700" swimtime="00:07:54.04" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1325" eventid="34" swimtime="00:04:13.67" lane="6" heatid="34005">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:58.35" />
                    <SPLIT distance="200" swimtime="00:02:05.09" />
                    <SPLIT distance="300" swimtime="00:03:11.25" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="366" birthdate="2006-01-01" gender="F" lastname="Jachmann" firstname="Valerie" license="0">
              <RESULTS>
                <RESULT resultid="1342" eventid="1" swimtime="00:00:20.12" lane="5" heatid="1013" />
                <RESULT resultid="1343" eventid="13" swimtime="00:00:40.11" lane="4" heatid="13006" />
                <RESULT resultid="1493" eventid="21" swimtime="00:00:39.38" lane="4" heatid="21001" />
                <RESULT resultid="1344" eventid="31" swimtime="00:00:45.80" lane="3" heatid="31017" />
                <RESULT resultid="1345" eventid="37" swimtime="00:00:18.03" lane="5" heatid="37006" />
                <RESULT resultid="1556" eventid="45" swimtime="00:00:18.15" lane="7" heatid="45001" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="367" birthdate="2003-01-01" gender="M" lastname="Schley" firstname="Wenzel" license="0">
              <RESULTS>
                <RESULT resultid="1346" eventid="10" swimtime="00:14:26.33" lane="3" heatid="10001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:49.62" />
                    <SPLIT distance="200" swimtime="00:01:44.72" />
                    <SPLIT distance="300" swimtime="00:02:41.86" />
                    <SPLIT distance="400" swimtime="00:03:39.98" />
                    <SPLIT distance="500" swimtime="00:04:38.35" />
                    <SPLIT distance="600" swimtime="00:05:36.64" />
                    <SPLIT distance="700" swimtime="00:06:35.52" />
                    <SPLIT distance="800" swimtime="00:07:34.28" />
                    <SPLIT distance="900" swimtime="00:08:33.12" />
                    <SPLIT distance="1000" swimtime="00:09:32.21" />
                    <SPLIT distance="1100" swimtime="00:10:31.33" />
                    <SPLIT distance="1200" swimtime="00:11:30.42" />
                    <SPLIT distance="1300" swimtime="00:12:29.35" />
                    <SPLIT distance="1400" swimtime="00:13:28.53" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1348" eventid="20" swimtime="00:03:23.46" lane="5" heatid="20002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:47.00" />
                    <SPLIT distance="200" swimtime="00:01:38.44" />
                    <SPLIT distance="300" swimtime="00:02:31.48" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1347" eventid="26" swimtime="00:07:19.57" lane="6" heatid="26001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:49.58" />
                    <SPLIT distance="200" swimtime="00:01:44.26" />
                    <SPLIT distance="300" swimtime="00:02:40.55" />
                    <SPLIT distance="400" swimtime="00:03:37.28" />
                    <SPLIT distance="500" swimtime="00:04:33.69" />
                    <SPLIT distance="600" swimtime="00:05:30.03" />
                    <SPLIT distance="700" swimtime="00:06:25.87" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1349" eventid="38" swimtime="00:00:17.15" lane="3" heatid="38008" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="368" birthdate="2008-01-01" gender="M" lastname="Stegemann" firstname="Wilhelm" license="0">
              <RESULTS>
                <RESULT resultid="1350" eventid="2" swimtime="00:00:18.95" lane="1" heatid="2009" />
                <RESULT resultid="1351" eventid="14" swimtime="00:00:43.23" lane="1" heatid="14005" />
                <RESULT resultid="1352" eventid="16" swimtime="00:01:39.17" lane="7" heatid="16006">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:48.57" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1353" eventid="32" swimtime="00:00:41.37" lane="4" heatid="32009" />
                <RESULT resultid="1354" eventid="38" swimtime="00:00:17.89" lane="7" heatid="38007" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY number="1" gender="M" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="1326" eventid="12" swimtime="00:06:39.09" lane="5" heatid="12002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:42.49" />
                    <SPLIT distance="200" swimtime="00:01:31.30" />
                    <SPLIT distance="300" swimtime="00:02:21.51" />
                    <SPLIT distance="400" swimtime="00:03:21.98" />
                    <SPLIT distance="500" swimtime="00:04:09.04" />
                    <SPLIT distance="600" swimtime="00:05:00.52" />
                    <SPLIT distance="700" swimtime="00:05:47.53" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="336" number="1" />
                    <RELAYPOSITION athleteid="335" number="2" />
                    <RELAYPOSITION athleteid="368" number="3" />
                    <RELAYPOSITION athleteid="367" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT resultid="1327" eventid="49" swimtime="00:02:47.20" lane="3" heatid="49002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:41.58" />
                    <SPLIT distance="200" swimtime="00:01:21.69" />
                    <SPLIT distance="300" swimtime="00:02:06.36" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="368" number="1" />
                    <RELAYPOSITION athleteid="336" number="2" />
                    <RELAYPOSITION athleteid="335" number="3" />
                    <RELAYPOSITION athleteid="367" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" gender="X" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="1328" eventid="30" swimtime="00:01:20.12" lane="5" heatid="30004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:40.05" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="367" number="1" />
                    <RELAYPOSITION athleteid="348" number="2" />
                    <RELAYPOSITION athleteid="337" number="3" />
                    <RELAYPOSITION athleteid="368" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" gender="F" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="1329" eventid="11" swimtime="00:07:07.82" lane="6" heatid="11003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:49.40" />
                    <SPLIT distance="200" swimtime="00:01:43.53" />
                    <SPLIT distance="300" swimtime="00:02:34.00" />
                    <SPLIT distance="400" swimtime="00:03:29.68" />
                    <SPLIT distance="500" swimtime="00:04:22.96" />
                    <SPLIT distance="600" swimtime="00:05:23.98" />
                    <SPLIT distance="700" swimtime="00:06:13.96" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="327" number="1" />
                    <RELAYPOSITION athleteid="348" number="2" />
                    <RELAYPOSITION athleteid="337" number="3" />
                    <RELAYPOSITION athleteid="366" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT resultid="1330" eventid="48" swimtime="00:03:05.81" lane="6" heatid="48003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:45.23" />
                    <SPLIT distance="200" swimtime="00:01:34.64" />
                    <SPLIT distance="300" swimtime="00:02:21.03" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="366" number="1" />
                    <RELAYPOSITION athleteid="333" number="2" />
                    <RELAYPOSITION athleteid="348" number="3" />
                    <RELAYPOSITION athleteid="327" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" gender="X" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="1331" eventid="30" status="DSQ" swimtime="00:01:15.75" lane="3" heatid="30004" comment="1. Schwimmer Falscher Start.">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:37.84" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="327" number="1" />
                    <RELAYPOSITION athleteid="336" number="2" />
                    <RELAYPOSITION athleteid="366" number="3" />
                    <RELAYPOSITION athleteid="335" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" gender="F" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="1332" eventid="11" swimtime="00:08:16.70" lane="8" heatid="11003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:57.88" />
                    <SPLIT distance="200" swimtime="00:02:01.48" />
                    <SPLIT distance="300" swimtime="00:03:05.38" />
                    <SPLIT distance="400" swimtime="00:04:12.96" />
                    <SPLIT distance="500" swimtime="00:05:11.72" />
                    <SPLIT distance="600" swimtime="00:06:17.92" />
                    <SPLIT distance="700" swimtime="00:07:13.62" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="333" number="1" />
                    <RELAYPOSITION athleteid="339" number="2" />
                    <RELAYPOSITION athleteid="341" number="3" />
                    <RELAYPOSITION athleteid="351" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" gender="F" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="1333" eventid="48" swimtime="00:03:36.52" lane="2" heatid="48003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:50.21" />
                    <SPLIT distance="200" swimtime="00:01:45.08" />
                    <SPLIT distance="300" swimtime="00:02:47.42" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="337" number="1" />
                    <RELAYPOSITION athleteid="341" number="2" />
                    <RELAYPOSITION athleteid="339" number="3" />
                    <RELAYPOSITION athleteid="351" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" gender="M" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="1334" eventid="12" swimtime="00:10:23.08" lane="4" heatid="12001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:02.62" />
                    <SPLIT distance="200" swimtime="00:02:09.23" />
                    <SPLIT distance="400" swimtime="00:05:13.14" />
                    <SPLIT distance="500" swimtime="00:06:30.68" />
                    <SPLIT distance="600" swimtime="00:07:51.11" />
                    <SPLIT distance="700" swimtime="00:09:04.34" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="347" number="1" />
                    <RELAYPOSITION athleteid="340" number="2" />
                    <RELAYPOSITION athleteid="331" number="3" />
                    <RELAYPOSITION athleteid="345" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT resultid="1335" eventid="49" swimtime="00:04:29.63" lane="3" heatid="49001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:16.71" />
                    <SPLIT distance="200" swimtime="00:02:23.70" />
                    <SPLIT distance="300" swimtime="00:03:24.37" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="331" number="1" />
                    <RELAYPOSITION athleteid="345" number="2" />
                    <RELAYPOSITION athleteid="347" number="3" />
                    <RELAYPOSITION athleteid="343" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" gender="F" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="1336" eventid="11" swimtime="00:09:31.18" lane="3" heatid="11001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:02.02" />
                    <SPLIT distance="200" swimtime="00:02:08.40" />
                    <SPLIT distance="300" swimtime="00:03:23.54" />
                    <SPLIT distance="400" swimtime="00:04:46.73" />
                    <SPLIT distance="500" swimtime="00:05:58.21" />
                    <SPLIT distance="600" swimtime="00:07:18.30" />
                    <SPLIT distance="700" swimtime="00:08:21.43" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="338" number="1" />
                    <RELAYPOSITION athleteid="342" number="2" />
                    <RELAYPOSITION athleteid="329" number="3" />
                    <RELAYPOSITION athleteid="344" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT resultid="1337" eventid="48" swimtime="00:04:17.23" lane="3" heatid="48001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:00.35" />
                    <SPLIT distance="200" swimtime="00:02:08.30" />
                    <SPLIT distance="300" swimtime="00:03:16.92" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="344" number="1" />
                    <RELAYPOSITION athleteid="342" number="2" />
                    <RELAYPOSITION athleteid="349" number="3" />
                    <RELAYPOSITION athleteid="338" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" gender="X" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="1338" eventid="30" swimtime="00:01:47.20" lane="4" heatid="30001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:52.41" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="347" number="1" />
                    <RELAYPOSITION athleteid="338" number="2" />
                    <RELAYPOSITION athleteid="352" number="3" />
                    <RELAYPOSITION athleteid="344" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" gender="F" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="1339" eventid="48" swimtime="00:04:36.69" lane="5" heatid="48001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:07.89" />
                    <SPLIT distance="200" swimtime="00:02:17.58" />
                    <SPLIT distance="300" swimtime="00:03:29.51" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="332" number="1" />
                    <RELAYPOSITION athleteid="330" number="2" />
                    <RELAYPOSITION athleteid="334" number="3" />
                    <RELAYPOSITION athleteid="329" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" gender="X" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="1340" eventid="30" swimtime="00:02:01.51" lane="5" heatid="30001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:00.68" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="349" number="1" />
                    <RELAYPOSITION athleteid="331" number="2" />
                    <RELAYPOSITION athleteid="329" number="3" />
                    <RELAYPOSITION athleteid="345" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" gender="X" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="1341" eventid="30" swimtime="00:01:53.36" lane="3" heatid="30001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:58.00" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="334" number="1" />
                    <RELAYPOSITION athleteid="343" number="2" />
                    <RELAYPOSITION athleteid="330" number="3" />
                    <RELAYPOSITION athleteid="353" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB name="TSC Schwandorf.de" nation="GER" region="34" code="0">
          <ATHLETES>
            <ATHLETE athleteid="68" birthdate="2007-01-01" gender="F" lastname="Rödl" firstname="Emily" license="0">
              <RESULTS>
                <RESULT resultid="228" eventid="9" swimtime="00:16:18.57" lane="1" heatid="9001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:59.47" />
                    <SPLIT distance="200" swimtime="00:02:04.20" />
                    <SPLIT distance="300" swimtime="00:03:10.43" />
                    <SPLIT distance="400" swimtime="00:04:17.23" />
                    <SPLIT distance="500" swimtime="00:05:23.77" />
                    <SPLIT distance="600" swimtime="00:06:30.80" />
                    <SPLIT distance="700" swimtime="00:07:36.94" />
                    <SPLIT distance="800" swimtime="00:08:43.41" />
                    <SPLIT distance="900" swimtime="00:09:49.84" />
                    <SPLIT distance="1000" swimtime="00:10:55.64" />
                    <SPLIT distance="1100" swimtime="00:12:02.04" />
                    <SPLIT distance="1200" swimtime="00:13:08.45" />
                    <SPLIT distance="1300" swimtime="00:14:14.64" />
                    <SPLIT distance="1400" swimtime="00:15:19.87" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="229" eventid="15" swimtime="00:01:48.47" lane="4" heatid="15009">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:52.37" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="230" eventid="17" swimtime="00:08:25.84" lane="6" heatid="17005">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:57.51" />
                    <SPLIT distance="200" swimtime="00:02:01.29" />
                    <SPLIT distance="300" swimtime="00:03:06.36" />
                    <SPLIT distance="400" swimtime="00:04:11.34" />
                    <SPLIT distance="500" swimtime="00:05:16.67" />
                    <SPLIT distance="600" swimtime="00:06:22.39" />
                    <SPLIT distance="700" swimtime="00:07:26.83" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="231" eventid="33" swimtime="00:03:59.04" lane="8" heatid="33007">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:55.45" />
                    <SPLIT distance="200" swimtime="00:01:57.16" />
                    <SPLIT distance="300" swimtime="00:03:00.00" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="232" eventid="37" swimtime="00:00:19.82" lane="6" heatid="37005" />
                <RESULT resultid="233" eventid="39" swimtime="00:00:25.53" lane="1" heatid="39004" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="69" birthdate="2011-01-01" gender="F" lastname="Maget" firstname="Matilda" license="0">
              <RESULTS>
                <RESULT resultid="234" eventid="1" swimtime="00:00:25.69" lane="7" heatid="1002" />
                <RESULT resultid="235" eventid="13" swimtime="00:01:09.98" lane="1" heatid="13001" />
                <RESULT resultid="236" eventid="15" swimtime="00:02:21.62" lane="6" heatid="15002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:08.71" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="237" eventid="31" swimtime="00:01:00.79" lane="8" heatid="31003" />
                <RESULT resultid="238" eventid="35" swimtime="00:00:26.69" lane="6" heatid="35001" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="70" birthdate="2010-01-01" gender="F" lastname="Seitz" firstname="Melina" license="0">
              <RESULTS>
                <RESULT resultid="239" eventid="1" swimtime="00:00:24.95" lane="5" heatid="1005" />
                <RESULT resultid="240" eventid="13" swimtime="00:00:57.71" lane="3" heatid="13002" />
                <RESULT resultid="241" eventid="15" swimtime="00:02:13.55" lane="6" heatid="15003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:05.50" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="242" eventid="31" swimtime="00:00:56.18" lane="1" heatid="31006" />
                <RESULT resultid="243" eventid="35" swimtime="00:00:25.38" lane="1" heatid="35002" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="71" birthdate="2004-01-01" gender="F" lastname="Kohler" firstname="Nina" license="0">
              <RESULTS>
                <RESULT resultid="244" eventid="1" swimtime="00:00:19.99" lane="3" heatid="1014" />
                <RESULT resultid="1410" eventid="7" swimtime="00:00:19.67" lane="8" heatid="7001" />
                <RESULT resultid="245" eventid="13" swimtime="00:00:40.72" lane="5" heatid="13006" />
                <RESULT resultid="246" eventid="15" swimtime="00:01:38.09" lane="5" heatid="15012">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:47.49" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1496" eventid="21" swimtime="00:00:40.99" lane="6" heatid="21001" />
                <RESULT resultid="1518" eventid="23" swimtime="00:01:40.38" lane="2" heatid="23001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:47.93" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="247" eventid="31" swimtime="00:00:43.77" lane="5" heatid="31015" />
                <RESULT resultid="248" eventid="37" swimtime="00:00:17.80" lane="3" heatid="37007" />
                <RESULT resultid="1540" eventid="41" swimtime="00:00:45.74" lane="7" heatid="41001" />
                <RESULT resultid="1553" eventid="45" swimtime="00:00:17.99" lane="3" heatid="45001" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="TSC Weimar e.V." nation="GER" region="35" code="174112">
          <ATHLETES>
            <ATHLETE athleteid="180" birthdate="2010-01-01" gender="F" lastname="Seyfarth" firstname="Annie" license="0">
              <RESULTS>
                <RESULT resultid="668" eventid="1" swimtime="00:00:27.97" lane="5" heatid="1002" />
                <RESULT resultid="669" eventid="15" swimtime="00:02:12.60" lane="3" heatid="15004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:01.91" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="670" eventid="31" swimtime="00:01:01.08" lane="2" heatid="31003" />
                <RESULT resultid="671" eventid="33" swimtime="00:04:46.20" lane="7" heatid="33002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:06.78" />
                    <SPLIT distance="200" swimtime="00:02:24.50" />
                    <SPLIT distance="300" swimtime="00:03:37.11" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="181" birthdate="2010-01-01" gender="M" lastname="Bellmann" firstname="Arvid" license="0">
              <RESULTS>
                <RESULT resultid="672" eventid="2" swimtime="00:00:25.71" lane="5" heatid="2003" />
                <RESULT resultid="673" eventid="14" swimtime="00:00:57.11" lane="3" heatid="14001" />
                <RESULT resultid="674" eventid="16" swimtime="00:02:12.85" lane="4" heatid="16002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:05.40" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="675" eventid="20" swimtime="00:05:08.64" lane="6" heatid="20001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:09.98" />
                    <SPLIT distance="200" swimtime="00:02:30.51" />
                    <SPLIT distance="300" swimtime="00:03:54.79" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="676" eventid="32" swimtime="00:00:57.90" lane="3" heatid="32003" />
                <RESULT resultid="677" eventid="34" swimtime="00:04:53.40" lane="8" heatid="34003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:08.31" />
                    <SPLIT distance="200" swimtime="00:02:23.99" />
                    <SPLIT distance="300" swimtime="00:03:44.24" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="678" eventid="36" swimtime="00:00:25.44" lane="3" heatid="36001" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="182" birthdate="2004-01-01" gender="M" lastname="Haufe" firstname="Elias" license="0">
              <RESULTS>
                <RESULT resultid="679" eventid="32" swimtime="00:00:44.93" lane="7" heatid="32009" />
                <RESULT resultid="680" eventid="38" swimtime="00:00:16.27" lane="5" heatid="38007" />
                <RESULT resultid="1564" eventid="46" swimtime="00:00:16.27" lane="7" heatid="46001" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="183" birthdate="2009-01-01" gender="M" lastname="Krebs" firstname="Emil" license="0">
              <RESULTS>
                <RESULT resultid="681" eventid="2" swimtime="00:00:25.46" lane="3" heatid="2002" />
                <RESULT resultid="682" eventid="38" swimtime="00:00:25.17" lane="1" heatid="38002" />
                <RESULT resultid="683" eventid="40" swimtime="00:00:26.07" lane="3" heatid="40002" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="184" birthdate="2007-01-01" gender="M" lastname="Röthlich" firstname="Finn" license="0">
              <RESULTS>
                <RESULT resultid="684" eventid="2" swimtime="00:00:22.33" lane="2" heatid="2007" />
                <RESULT resultid="688" eventid="6" swimtime="00:00:53.00" lane="5" heatid="6003" />
                <RESULT resultid="685" eventid="14" swimtime="00:00:50.64" lane="1" heatid="14003" />
                <RESULT resultid="686" eventid="32" swimtime="00:00:52.23" lane="4" heatid="32005" />
                <RESULT resultid="687" eventid="38" swimtime="00:00:20.21" lane="6" heatid="38005" />
                <RESULT resultid="689" eventid="40" swimtime="00:00:23.43" lane="3" heatid="40003" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="185" birthdate="2005-01-01" gender="M" lastname="Linne" firstname="Georg" license="0">
              <RESULTS>
                <RESULT resultid="690" eventid="14" swimtime="00:00:39.36" lane="5" heatid="14004" />
                <RESULT resultid="691" eventid="16" swimtime="00:01:35.34" lane="2" heatid="16007">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:45.21" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1510" eventid="22" swimtime="00:00:39.40" lane="1" heatid="22001" />
                <RESULT resultid="1532" eventid="24" swimtime="00:01:38.10" lane="7" heatid="24001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:46.38" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="692" eventid="28" swimtime="00:03:14.63" lane="3" heatid="28001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:44.75" />
                    <SPLIT distance="200" swimtime="00:01:34.28" />
                    <SPLIT distance="300" swimtime="00:02:25.86" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="693" eventid="32" swimtime="00:00:43.61" lane="6" heatid="32009" />
                <RESULT resultid="694" eventid="34" swimtime="00:03:30.49" lane="4" heatid="34006">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:47.53" />
                    <SPLIT distance="200" swimtime="00:01:40.57" />
                    <SPLIT distance="300" swimtime="00:02:35.72" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="695" eventid="38" swimtime="00:00:17.54" lane="7" heatid="38009" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="186" birthdate="2009-01-01" gender="M" lastname="Klabunde" firstname="Kalle" license="0">
              <RESULTS>
                <RESULT resultid="696" eventid="34" swimtime="00:04:46.77" lane="5" heatid="34002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:04.24" />
                    <SPLIT distance="200" swimtime="00:02:16.28" />
                    <SPLIT distance="300" swimtime="00:03:25.03" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="697" eventid="38" swimtime="00:00:26.50" lane="7" heatid="38002" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="187" birthdate="2010-01-01" gender="F" lastname="Pontes" firstname="Lena" license="0">
              <RESULTS>
                <RESULT resultid="698" eventid="1" swimtime="00:00:26.98" lane="3" heatid="1004" />
                <RESULT resultid="699" eventid="31" swimtime="00:00:58.68" lane="8" heatid="31004" />
                <RESULT resultid="700" eventid="35" swimtime="00:00:25.78" lane="7" heatid="35002" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="188" birthdate="2011-01-01" gender="M" lastname="Bellmann" firstname="Lennart" license="0">
              <RESULTS>
                <RESULT resultid="701" eventid="2" swimtime="00:00:24.36" lane="4" heatid="2004" />
                <RESULT resultid="702" eventid="14" swimtime="00:01:01.17" lane="7" heatid="14001" />
                <RESULT resultid="703" eventid="16" swimtime="00:02:04.31" lane="4" heatid="16003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:59.69" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="704" eventid="32" swimtime="00:00:55.14" lane="8" heatid="32005" />
                <RESULT resultid="705" eventid="34" swimtime="00:04:27.04" lane="1" heatid="34004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:03.95" />
                    <SPLIT distance="200" swimtime="00:02:12.10" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="706" eventid="36" swimtime="00:00:25.28" lane="6" heatid="36001" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="189" birthdate="2011-01-01" gender="F" lastname="Hüttig" firstname="Maline" license="0">
              <RESULTS>
                <RESULT resultid="707" eventid="1" swimtime="00:00:29.51" lane="8" heatid="1003" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="190" birthdate="1971-01-01" gender="F" lastname="Klabunde" firstname="Monique" license="0">
              <RESULTS>
                <RESULT resultid="708" eventid="15" swimtime="00:01:59.62" lane="6" heatid="15006">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:57.30" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="709" eventid="31" swimtime="00:00:54.17" lane="6" heatid="31009" />
                <RESULT resultid="710" eventid="33" swimtime="00:04:17.84" lane="7" heatid="33005">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:59.35" />
                    <SPLIT distance="200" swimtime="00:02:04.82" />
                    <SPLIT distance="300" swimtime="00:03:11.88" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="191" birthdate="2004-01-01" gender="M" lastname="Röthlich" firstname="Nils" license="0">
              <RESULTS>
                <RESULT resultid="711" eventid="14" swimtime="00:00:46.77" lane="4" heatid="14003" />
                <RESULT resultid="712" eventid="32" swimtime="00:00:48.18" lane="2" heatid="32008" />
                <RESULT resultid="713" eventid="38" swimtime="00:00:19.96" lane="7" heatid="38006" />
                <RESULT resultid="714" eventid="40" swimtime="00:00:24.83" lane="7" heatid="40003" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="192" birthdate="2008-01-01" gender="M" lastname="Kraft" firstname="Simon" license="0">
              <RESULTS>
                <RESULT resultid="715" eventid="2" swimtime="00:00:20.07" lane="2" heatid="2008" />
                <RESULT resultid="716" eventid="14" swimtime="00:00:40.96" lane="6" heatid="14004" />
                <RESULT resultid="717" eventid="20" status="DNS" swimtime="00:00:00.00" lane="7" heatid="20002" />
                <RESULT resultid="1502" eventid="22" status="WDR" swimtime="00:00:00.00" lane="0" heatid="22000" />
                <RESULT resultid="718" eventid="32" swimtime="00:00:44.39" lane="7" heatid="32008" />
                <RESULT resultid="719" eventid="38" swimtime="00:00:17.62" lane="8" heatid="38009" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="193" birthdate="2006-01-01" gender="M" lastname="Hauser" firstname="Theo" license="0">
              <RESULTS>
                <RESULT resultid="720" eventid="2" swimtime="00:00:20.20" lane="4" heatid="2008" />
                <RESULT resultid="721" eventid="14" swimtime="00:00:45.36" lane="5" heatid="14003" />
                <RESULT resultid="722" eventid="32" swimtime="00:00:45.44" lane="8" heatid="32009" />
                <RESULT resultid="723" eventid="38" swimtime="00:00:18.93" lane="8" heatid="38007" />
                <RESULT resultid="724" eventid="40" swimtime="00:00:22.45" lane="6" heatid="40004" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY number="1" gender="M" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="664" eventid="49" swimtime="00:03:54.72" lane="8" heatid="49002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:50.90" />
                    <SPLIT distance="200" swimtime="00:01:52.30" />
                    <SPLIT distance="300" swimtime="00:02:54.18" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="192" number="1" />
                    <RELAYPOSITION athleteid="186" number="2" />
                    <RELAYPOSITION athleteid="183" number="3" />
                    <RELAYPOSITION athleteid="181" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="2" gender="X" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="665" eventid="30" swimtime="00:01:38.90" lane="2" heatid="30002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:46.77" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="192" number="1" />
                    <RELAYPOSITION athleteid="187" number="2" />
                    <RELAYPOSITION athleteid="180" number="3" />
                    <RELAYPOSITION athleteid="181" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="3" gender="M" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="666" eventid="49" swimtime="00:02:57.98" lane="2" heatid="49002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:45.14" />
                    <SPLIT distance="200" swimtime="00:01:29.11" />
                    <SPLIT distance="300" swimtime="00:02:15.89" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="182" number="1" />
                    <RELAYPOSITION athleteid="193" number="2" />
                    <RELAYPOSITION athleteid="191" number="3" />
                    <RELAYPOSITION athleteid="185" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="4" gender="M" agemin="-1" agemax="-1" agetotalmin="-1" agetotalmax="-1" name="">
              <RESULTS>
                <RESULT resultid="667" eventid="12" swimtime="00:08:30.68" lane="8" heatid="12002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:55.62" />
                    <SPLIT distance="200" swimtime="00:01:56.44" />
                    <SPLIT distance="300" swimtime="00:02:56.56" />
                    <SPLIT distance="400" swimtime="00:04:02.49" />
                    <SPLIT distance="500" swimtime="00:05:09.84" />
                    <SPLIT distance="600" swimtime="00:06:19.31" />
                    <SPLIT distance="700" swimtime="00:07:18.59" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="192" number="1" />
                    <RELAYPOSITION athleteid="193" number="2" />
                    <RELAYPOSITION athleteid="181" number="3" />
                    <RELAYPOSITION athleteid="184" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB name="TSG Schwäbisch Hall" nation="GER" region="18" code="2545">
          <ATHLETES>
            <ATHLETE athleteid="130" birthdate="1967-01-01" gender="M" lastname="Lochstampfer" firstname="Gunter" license="78798">
              <RESULTS>
                <RESULT resultid="479" eventid="2" swimtime="00:00:23.87" lane="6" heatid="2005" />
                <RESULT resultid="482" eventid="6" swimtime="00:00:54.45" lane="3" heatid="6003" />
                <RESULT resultid="480" eventid="32" swimtime="00:00:54.02" lane="5" heatid="32005" />
                <RESULT resultid="481" eventid="38" swimtime="00:00:22.37" lane="8" heatid="38002" />
                <RESULT resultid="483" eventid="40" swimtime="00:00:25.30" lane="1" heatid="40003" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="TSG TU Ilmenau 56 e.V." nation="GER" region="35" code="0">
          <ATHLETES>
            <ATHLETE athleteid="369" birthdate="2009-01-01" gender="F" lastname="Weber" firstname="Augusta Swantje" license="0">
              <RESULTS>
                <RESULT resultid="1355" eventid="1" swimtime="00:00:27.42" lane="4" heatid="1003" />
                <RESULT resultid="1356" eventid="13" swimtime="00:01:05.21" lane="5" heatid="13001" />
                <RESULT resultid="1357" eventid="15" swimtime="00:02:20.49" lane="3" heatid="15003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:07.16" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1358" eventid="31" swimtime="00:01:02.87" lane="1" heatid="31004" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="370" birthdate="2001-01-01" gender="M" lastname="Pohl" firstname="Enrico" license="0">
              <RESULTS>
                <RESULT resultid="1359" eventid="14" swimtime="00:00:38.50" lane="3" heatid="14006" />
                <RESULT resultid="1360" eventid="16" swimtime="00:01:34.26" lane="6" heatid="16008">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:44.07" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1509" eventid="22" swimtime="00:00:37.02" lane="7" heatid="22001" />
                <RESULT resultid="1526" eventid="24" status="WDR" swimtime="00:00:00.00" lane="0" heatid="24000" />
                <RESULT resultid="1361" eventid="32" swimtime="00:00:39.09" lane="5" heatid="32011" />
                <RESULT resultid="1362" eventid="38" swimtime="00:00:15.95" lane="5" heatid="38008" />
                <RESULT resultid="1546" eventid="42" swimtime="00:00:38.19" lane="6" heatid="42001" />
                <RESULT resultid="1563" eventid="46" swimtime="00:00:15.84" lane="2" heatid="46001" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="371" birthdate="2008-01-01" gender="F" lastname="Liebhold" firstname="Lotta" license="0">
              <RESULTS>
                <RESULT resultid="1363" eventid="1" swimtime="00:00:25.80" lane="8" heatid="1007" />
                <RESULT resultid="1364" eventid="15" swimtime="00:02:08.49" lane="4" heatid="15005">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:01.35" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1365" eventid="17" swimtime="00:09:35.00" lane="7" heatid="17003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:03.61" />
                    <SPLIT distance="200" swimtime="00:02:15.94" />
                    <SPLIT distance="300" swimtime="00:03:30.36" />
                    <SPLIT distance="400" swimtime="00:04:45.28" />
                    <SPLIT distance="500" swimtime="00:06:00.92" />
                    <SPLIT distance="600" swimtime="00:07:16.18" />
                    <SPLIT distance="700" swimtime="00:08:28.77" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1366" eventid="31" swimtime="00:00:57.04" lane="8" heatid="31008" />
                <RESULT resultid="1367" eventid="33" swimtime="00:04:29.02" lane="3" heatid="33003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:00.45" />
                    <SPLIT distance="200" swimtime="00:02:10.36" />
                    <SPLIT distance="300" swimtime="00:03:22.05" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="372" birthdate="2007-01-01" gender="M" lastname="Stuwe" firstname="Paul" license="0">
              <RESULTS>
                <RESULT resultid="1368" eventid="2" swimtime="00:00:22.99" lane="3" heatid="2006" />
                <RESULT resultid="1369" eventid="4" swimtime="00:19:56.16" lane="4" heatid="4001">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:06.36" />
                    <SPLIT distance="200" swimtime="00:02:21.55" />
                    <SPLIT distance="300" swimtime="00:03:38.68" />
                    <SPLIT distance="400" swimtime="00:04:57.85" />
                    <SPLIT distance="500" swimtime="00:06:17.67" />
                    <SPLIT distance="600" swimtime="00:07:38.37" />
                    <SPLIT distance="700" swimtime="00:08:59.95" />
                    <SPLIT distance="800" swimtime="00:10:23.04" />
                    <SPLIT distance="900" swimtime="00:11:45.85" />
                    <SPLIT distance="1000" swimtime="00:13:06.93" />
                    <SPLIT distance="1100" swimtime="00:14:28.59" />
                    <SPLIT distance="1200" swimtime="00:15:50.77" />
                    <SPLIT distance="1300" swimtime="00:17:13.34" />
                    <SPLIT distance="1400" swimtime="00:18:34.86" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1370" eventid="14" swimtime="00:00:48.49" lane="2" heatid="14003" />
                <RESULT resultid="1371" eventid="18" swimtime="00:09:07.89" lane="2" heatid="18003">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:00.66" />
                    <SPLIT distance="200" swimtime="00:02:07.17" />
                    <SPLIT distance="300" swimtime="00:03:16.29" />
                    <SPLIT distance="400" swimtime="00:04:26.74" />
                    <SPLIT distance="500" swimtime="00:05:38.69" />
                    <SPLIT distance="600" swimtime="00:06:50.06" />
                    <SPLIT distance="700" swimtime="00:07:59.74" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1372" eventid="20" swimtime="00:04:20.37" lane="2" heatid="20002">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:57.50" />
                    <SPLIT distance="200" swimtime="00:02:04.41" />
                    <SPLIT distance="300" swimtime="00:03:13.38" />
                  </SPLITS>
                </RESULT>
                <RESULT resultid="1373" eventid="32" swimtime="00:00:50.84" lane="4" heatid="32006" />
                <RESULT resultid="1374" eventid="34" swimtime="00:04:12.04" lane="7" heatid="34004">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:57.03" />
                    <SPLIT distance="200" swimtime="00:02:00.05" />
                    <SPLIT distance="300" swimtime="00:03:06.63" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
      </CLUBS>
    </MEET>
  </MEETS>
  <TIMESTANDARDLISTS>
    <TIMESTANDARDLIST name="Pflichtzeiten 1958 und jünger weiblich" course="LCM" gender="F" timestandardlistid="1">
      <AGEGROUP agemax="-1" agemin="65" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:07:00.00">
          <SWIMSTYLE distance="400" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:13:00.00">
          <SWIMSTYLE distance="800" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:39.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="APNEA" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:35.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:06:55.00">
          <SWIMSTYLE distance="400" relaycount="1" stroke="IMMERSION" technique="DIVE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:20.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:34.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="IMMERSION" technique="DIVE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:07:00.00">
          <SWIMSTYLE distance="400" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:17:50.00">
          <SWIMSTYLE distance="1500" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:17:50.00">
          <SWIMSTYLE distance="1500" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:13:00.00">
          <SWIMSTYLE distance="800" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:06:55.00">
          <SWIMSTYLE distance="400" relaycount="1" stroke="IMMERSION" technique="DIVE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:40.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST name="Pflichtzeiten 1959 bis 1969 weiblich" course="LCM" gender="F" timestandardlistid="2">
      <AGEGROUP agemax="64" agemin="54" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:06:20.00">
          <SWIMSTYLE distance="400" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:12:00.00">
          <SWIMSTYLE distance="800" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:35.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="APNEA" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:25.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:06:15.00">
          <SWIMSTYLE distance="400" relaycount="1" stroke="IMMERSION" technique="DIVE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:00.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:24.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="IMMERSION" technique="DIVE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:06:20.00">
          <SWIMSTYLE distance="400" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:12:00.00">
          <SWIMSTYLE distance="800" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:06:15.00">
          <SWIMSTYLE distance="400" relaycount="1" stroke="IMMERSION" technique="DIVE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:36.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST name="Pflichtzeiten 1969 bis 1978 weiblich" course="LCM" gender="F" timestandardlistid="3">
      <AGEGROUP agemax="54" agemin="45" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:05:20.00">
          <SWIMSTYLE distance="400" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:15.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:05:15.00">
          <SWIMSTYLE distance="400" relaycount="1" stroke="IMMERSION" technique="DIVE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:40.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:14.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="IMMERSION" technique="DIVE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:11:15.00">
          <SWIMSTYLE distance="800" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:31.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="APNEA" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:05:20.00">
          <SWIMSTYLE distance="400" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:17:50.00">
          <SWIMSTYLE distance="1500" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:17:50.00">
          <SWIMSTYLE distance="1500" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:11:15.00">
          <SWIMSTYLE distance="800" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:05:15.00">
          <SWIMSTYLE distance="400" relaycount="1" stroke="IMMERSION" technique="DIVE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:32.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST name="Pflichtzeiten 1979 bis 1988 weiblich" course="LCM" gender="F" timestandardlistid="4">
      <AGEGROUP agemax="44" agemin="35" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:04:55.00">
          <SWIMSTYLE distance="400" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:06.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:04:50.00">
          <SWIMSTYLE distance="400" relaycount="1" stroke="IMMERSION" technique="DIVE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:25.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:00.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="IMMERSION" technique="DIVE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:10:30.00">
          <SWIMSTYLE distance="800" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:28.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="APNEA" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:04:55.00">
          <SWIMSTYLE distance="400" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:17:50.00">
          <SWIMSTYLE distance="1500" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:17:50.00">
          <SWIMSTYLE distance="1500" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:10:30.00">
          <SWIMSTYLE distance="800" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:04:50.00">
          <SWIMSTYLE distance="400" relaycount="1" stroke="IMMERSION" technique="DIVE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:29.90">
          <SWIMSTYLE distance="50" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST name="Pflichtzeiten 1989 bis 1994 weiblich" course="LCM" gender="F" timestandardlistid="5">
      <AGEGROUP agemax="34" agemin="29" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:04:45.00">
          <SWIMSTYLE distance="400" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:01.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:04:40.00">
          <SWIMSTYLE distance="400" relaycount="1" stroke="IMMERSION" technique="DIVE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:10.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:00.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="IMMERSION" technique="DIVE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:10:00.00">
          <SWIMSTYLE distance="800" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:27.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="APNEA" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:04:45.00">
          <SWIMSTYLE distance="400" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:17:50.00">
          <SWIMSTYLE distance="1500" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:17:50.00">
          <SWIMSTYLE distance="1500" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:10:00.00">
          <SWIMSTYLE distance="800" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:04:40.00">
          <SWIMSTYLE distance="400" relaycount="1" stroke="IMMERSION" technique="DIVE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:28.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST name="Pflichtzeiten 1995 bis 2001 weiblich" course="LCM" gender="F" timestandardlistid="6">
      <AGEGROUP agemax="28" agemin="22" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:04:20.00">
          <SWIMSTYLE distance="400" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:54.50">
          <SWIMSTYLE distance="100" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:04:15.00">
          <SWIMSTYLE distance="400" relaycount="1" stroke="IMMERSION" technique="DIVE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:00.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:53.50">
          <SWIMSTYLE distance="100" relaycount="1" stroke="IMMERSION" technique="DIVE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:09:10.00">
          <SWIMSTYLE distance="800" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:22.50">
          <SWIMSTYLE distance="50" relaycount="1" stroke="APNEA" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:04:20.00">
          <SWIMSTYLE distance="400" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:17:50.00">
          <SWIMSTYLE distance="1500" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:17:50.00">
          <SWIMSTYLE distance="1500" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:09:10.00">
          <SWIMSTYLE distance="800" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:04:15.00">
          <SWIMSTYLE distance="400" relaycount="1" stroke="IMMERSION" technique="DIVE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:24.50">
          <SWIMSTYLE distance="50" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST name="Pflichtzeiten 2002 bis 2005 weiblich" course="LCM" gender="F" timestandardlistid="7">
      <AGEGROUP agemax="21" agemin="18" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:04:24.00">
          <SWIMSTYLE distance="400" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:54.50">
          <SWIMSTYLE distance="100" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:04:19.00">
          <SWIMSTYLE distance="400" relaycount="1" stroke="IMMERSION" technique="DIVE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:01.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:53.50">
          <SWIMSTYLE distance="100" relaycount="1" stroke="IMMERSION" technique="DIVE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:09:18.00">
          <SWIMSTYLE distance="800" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:22.50">
          <SWIMSTYLE distance="50" relaycount="1" stroke="APNEA" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:04:24.00">
          <SWIMSTYLE distance="400" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:18:07.00">
          <SWIMSTYLE distance="1500" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:18:07.00">
          <SWIMSTYLE distance="1500" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:09:18.00">
          <SWIMSTYLE distance="800" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:04:19.00">
          <SWIMSTYLE distance="400" relaycount="1" stroke="IMMERSION" technique="DIVE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:24.50">
          <SWIMSTYLE distance="50" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST name="Pflichtzeiten 2006 weiblich" course="LCM" gender="F" timestandardlistid="8">
      <AGEGROUP agemax="17" agemin="17" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:04:40.00">
          <SWIMSTYLE distance="400" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:58.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:04:40.00">
          <SWIMSTYLE distance="400" relaycount="1" stroke="IMMERSION" technique="DIVE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:08.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:58.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="IMMERSION" technique="DIVE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:09:53.00">
          <SWIMSTYLE distance="800" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:23.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="APNEA" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:04:40.00">
          <SWIMSTYLE distance="400" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:19:17.00">
          <SWIMSTYLE distance="1500" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:19:17.00">
          <SWIMSTYLE distance="1500" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:09:53.00">
          <SWIMSTYLE distance="800" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:04:40.00">
          <SWIMSTYLE distance="400" relaycount="1" stroke="IMMERSION" technique="DIVE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:25.80">
          <SWIMSTYLE distance="50" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST name="Pflichtzeiten 2007 weiblich" course="LCM" gender="F" timestandardlistid="9">
      <AGEGROUP agemax="16" agemin="16" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:04:45.00">
          <SWIMSTYLE distance="400" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:59.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:04:50.00">
          <SWIMSTYLE distance="400" relaycount="1" stroke="IMMERSION" technique="DIVE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:10.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:00.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="IMMERSION" technique="DIVE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:10:04.00">
          <SWIMSTYLE distance="800" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:23.50">
          <SWIMSTYLE distance="50" relaycount="1" stroke="APNEA" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:04:45.00">
          <SWIMSTYLE distance="400" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:19:37.00">
          <SWIMSTYLE distance="1500" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:19:37.00">
          <SWIMSTYLE distance="1500" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:10:04.00">
          <SWIMSTYLE distance="800" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:04:50.00">
          <SWIMSTYLE distance="400" relaycount="1" stroke="IMMERSION" technique="DIVE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:26.30">
          <SWIMSTYLE distance="50" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST name="Pflichtzeiten 2008 weiblich" course="LCM" gender="F" timestandardlistid="10">
      <AGEGROUP agemax="15" agemin="15" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:04:50.00">
          <SWIMSTYLE distance="400" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:00.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:05:00.00">
          <SWIMSTYLE distance="400" relaycount="1" stroke="IMMERSION" technique="DIVE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:13.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:02.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="IMMERSION" technique="DIVE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:10:14.00">
          <SWIMSTYLE distance="800" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:24.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="APNEA" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:04:50.00">
          <SWIMSTYLE distance="400" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:19:57.00">
          <SWIMSTYLE distance="1500" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:19:57.00">
          <SWIMSTYLE distance="1500" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:10:14.00">
          <SWIMSTYLE distance="800" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:05:00.00">
          <SWIMSTYLE distance="400" relaycount="1" stroke="IMMERSION" technique="DIVE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:26.70">
          <SWIMSTYLE distance="50" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST name="Pflichtzeiten 2009 weiblich" course="LCM" gender="F" timestandardlistid="11">
      <AGEGROUP agemax="14" agemin="14" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:05:00.00">
          <SWIMSTYLE distance="400" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:02.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:05:09.00">
          <SWIMSTYLE distance="400" relaycount="1" stroke="IMMERSION" technique="DIVE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:17.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:04.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="IMMERSION" technique="DIVE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:10:34.00">
          <SWIMSTYLE distance="800" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:25.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="APNEA" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:05:00.00">
          <SWIMSTYLE distance="400" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:20:36.00">
          <SWIMSTYLE distance="1500" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:20:36.00">
          <SWIMSTYLE distance="1500" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:10:34.00">
          <SWIMSTYLE distance="800" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:05:09.00">
          <SWIMSTYLE distance="400" relaycount="1" stroke="IMMERSION" technique="DIVE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:27.50">
          <SWIMSTYLE distance="50" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST name="Pflichtzeiten 2010 weiblich" course="LCM" gender="F" timestandardlistid="12">
      <AGEGROUP agemax="13" agemin="13" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:05:10.00">
          <SWIMSTYLE distance="400" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:27.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="IMMERSION" technique="DIVE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:05.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:05:30.00">
          <SWIMSTYLE distance="400" relaycount="1" stroke="IMMERSION" technique="DIVE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:24.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:10:50.00">
          <SWIMSTYLE distance="800" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:05:10.00">
          <SWIMSTYLE distance="400" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:06.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="IMMERSION" technique="DIVE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:20:56.00">
          <SWIMSTYLE distance="1500" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:20:56.00">
          <SWIMSTYLE distance="1500" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:10:50.00">
          <SWIMSTYLE distance="800" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:05:30.00">
          <SWIMSTYLE distance="400" relaycount="1" stroke="IMMERSION" technique="DIVE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:29.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST name="Pflichtzeiten 2011 weiblich" course="LCM" gender="F" timestandardlistid="13">
      <AGEGROUP agemax="12" agemin="12" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:05:25.00">
          <SWIMSTYLE distance="400" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:28.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="IMMERSION" technique="DIVE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:08.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:05:55.00">
          <SWIMSTYLE distance="400" relaycount="1" stroke="IMMERSION" technique="DIVE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:30.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:11:20.00">
          <SWIMSTYLE distance="800" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:05:25.00">
          <SWIMSTYLE distance="400" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:10.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="IMMERSION" technique="DIVE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:21:26.00">
          <SWIMSTYLE distance="1500" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:21:26.00">
          <SWIMSTYLE distance="1500" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:11:20.00">
          <SWIMSTYLE distance="800" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:05:55.00">
          <SWIMSTYLE distance="400" relaycount="1" stroke="IMMERSION" technique="DIVE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:30.50">
          <SWIMSTYLE distance="50" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST name="Pflichtzeiten 1958 und jünger männlich" course="LCM" gender="M" timestandardlistid="14">
      <AGEGROUP agemax="-1" agemin="65" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:06:40.00">
          <SWIMSTYLE distance="400" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:22.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:17:10.00">
          <SWIMSTYLE distance="1500" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:06:35.00">
          <SWIMSTYLE distance="400" relaycount="1" stroke="IMMERSION" technique="DIVE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:31.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="APNEA" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:12:30.00">
          <SWIMSTYLE distance="800" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:06:40.00">
          <SWIMSTYLE distance="400" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:17:10.00">
          <SWIMSTYLE distance="1500" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:33.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:19.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="IMMERSION" technique="DIVE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:12:30.00">
          <SWIMSTYLE distance="800" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:06:35.00">
          <SWIMSTYLE distance="400" relaycount="1" stroke="IMMERSION" technique="DIVE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:10.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST name="Pflichtzeiten 1959 bis 1969 männlich" course="LCM" gender="M" timestandardlistid="15">
      <AGEGROUP agemax="64" agemin="54" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:05:40.00">
          <SWIMSTYLE distance="400" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:10.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:05:40.00">
          <SWIMSTYLE distance="400" relaycount="1" stroke="IMMERSION" technique="DIVE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:28.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="APNEA" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:11:30.00">
          <SWIMSTYLE distance="800" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:05:40.00">
          <SWIMSTYLE distance="400" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:30.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:07.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="IMMERSION" technique="DIVE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:11:30.00">
          <SWIMSTYLE distance="800" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:05:40.00">
          <SWIMSTYLE distance="400" relaycount="1" stroke="IMMERSION" technique="DIVE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:40.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST name="Pflichtzeiten 1969 bis 1978 männlich" course="LCM" gender="M" timestandardlistid="16">
      <AGEGROUP agemax="54" agemin="45" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:05:10.00">
          <SWIMSTYLE distance="400" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:17:10.00">
          <SWIMSTYLE distance="1500" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:06.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:17:10.00">
          <SWIMSTYLE distance="1500" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:26.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="APNEA" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:10:45.00">
          <SWIMSTYLE distance="800" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:05:10.00">
          <SWIMSTYLE distance="400" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:05:05.00">
          <SWIMSTYLE distance="400" relaycount="1" stroke="IMMERSION" technique="DIVE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:28.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:03.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="IMMERSION" technique="DIVE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:10:45.00">
          <SWIMSTYLE distance="800" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:05:05.00">
          <SWIMSTYLE distance="400" relaycount="1" stroke="IMMERSION" technique="DIVE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:20.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST name="Pflichtzeiten 1979 bis 1988 männlich" course="LCM" gender="M" timestandardlistid="17">
      <AGEGROUP agemax="44" agemin="35" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:04:45.00">
          <SWIMSTYLE distance="400" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:17:10.00">
          <SWIMSTYLE distance="1500" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:58.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:17:10.00">
          <SWIMSTYLE distance="1500" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:23.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="APNEA" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:10:00.00">
          <SWIMSTYLE distance="800" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:04:45.00">
          <SWIMSTYLE distance="400" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:04:40.00">
          <SWIMSTYLE distance="400" relaycount="1" stroke="IMMERSION" technique="DIVE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:26.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:55.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="IMMERSION" technique="DIVE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:10:00.00">
          <SWIMSTYLE distance="800" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:04:40.00">
          <SWIMSTYLE distance="400" relaycount="1" stroke="IMMERSION" technique="DIVE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:10.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST name="Pflichtzeiten 1989 bis 1994 männlich" course="LCM" gender="M" timestandardlistid="18">
      <AGEGROUP agemax="34" agemin="29" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:04:20.00">
          <SWIMSTYLE distance="400" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:17:10.00">
          <SWIMSTYLE distance="1500" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:56.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:17:10.00">
          <SWIMSTYLE distance="1500" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:22.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="APNEA" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:09:30.00">
          <SWIMSTYLE distance="800" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:04:20.00">
          <SWIMSTYLE distance="400" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:04:15.00">
          <SWIMSTYLE distance="400" relaycount="1" stroke="IMMERSION" technique="DIVE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:25.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:53.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="IMMERSION" technique="DIVE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:09:30.00">
          <SWIMSTYLE distance="800" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:04:15.00">
          <SWIMSTYLE distance="400" relaycount="1" stroke="IMMERSION" technique="DIVE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:00.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST name="Pflichtzeiten 1995 bis 2001 männlich" course="LCM" gender="M" timestandardlistid="19">
      <AGEGROUP agemax="28" agemin="22" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:04:05.00">
          <SWIMSTYLE distance="400" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:17:10.00">
          <SWIMSTYLE distance="1500" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:51.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:17:10.00">
          <SWIMSTYLE distance="1500" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:20.50">
          <SWIMSTYLE distance="50" relaycount="1" stroke="APNEA" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:08:05.00">
          <SWIMSTYLE distance="800" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:04:05.00">
          <SWIMSTYLE distance="400" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:57.00">
          <SWIMSTYLE distance="400" relaycount="1" stroke="IMMERSION" technique="DIVE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:23.50">
          <SWIMSTYLE distance="50" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:49.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="IMMERSION" technique="DIVE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:08:05.00">
          <SWIMSTYLE distance="800" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:57.00">
          <SWIMSTYLE distance="400" relaycount="1" stroke="IMMERSION" technique="DIVE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:55.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST name="Pflichtzeiten 2002 bis 2005 männlich" course="LCM" gender="M" timestandardlistid="20">
      <AGEGROUP agemax="21" agemin="18" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:04:14.00">
          <SWIMSTYLE distance="400" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:17:27.00">
          <SWIMSTYLE distance="1500" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:52.20">
          <SWIMSTYLE distance="100" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:17:27.00">
          <SWIMSTYLE distance="1500" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:20.50">
          <SWIMSTYLE distance="50" relaycount="1" stroke="APNEA" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:08:57.00">
          <SWIMSTYLE distance="800" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:04:14.00">
          <SWIMSTYLE distance="400" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:57.00">
          <SWIMSTYLE distance="400" relaycount="1" stroke="IMMERSION" technique="DIVE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:24.50">
          <SWIMSTYLE distance="50" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:49.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="IMMERSION" technique="DIVE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:08:57.00">
          <SWIMSTYLE distance="800" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:57.00">
          <SWIMSTYLE distance="400" relaycount="1" stroke="IMMERSION" technique="DIVE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:57.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST name="Pflichtzeiten 2006 männlich" course="LCM" gender="M" timestandardlistid="21">
      <AGEGROUP agemax="17" agemin="17" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:04:35.00">
          <SWIMSTYLE distance="400" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:18:57.00">
          <SWIMSTYLE distance="1500" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:57.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:18:57.00">
          <SWIMSTYLE distance="1500" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:21.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="APNEA" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:09:43.00">
          <SWIMSTYLE distance="800" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:04:35.00">
          <SWIMSTYLE distance="400" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:04:26.00">
          <SWIMSTYLE distance="400" relaycount="1" stroke="IMMERSION" technique="DIVE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:25.40">
          <SWIMSTYLE distance="50" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:55.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="IMMERSION" technique="DIVE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:09:43.00">
          <SWIMSTYLE distance="800" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:04:26.00">
          <SWIMSTYLE distance="400" relaycount="1" stroke="IMMERSION" technique="DIVE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:06.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST name="Pflichtzeiten 2007 männlich" course="LCM" gender="M" timestandardlistid="22">
      <AGEGROUP agemax="16" agemin="16" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:04:40.00">
          <SWIMSTYLE distance="400" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:19:17.00">
          <SWIMSTYLE distance="1500" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:58.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:19:17.00">
          <SWIMSTYLE distance="1500" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:21.50">
          <SWIMSTYLE distance="50" relaycount="1" stroke="APNEA" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:09:53.00">
          <SWIMSTYLE distance="800" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:04:40.00">
          <SWIMSTYLE distance="400" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:04:40.00">
          <SWIMSTYLE distance="400" relaycount="1" stroke="IMMERSION" technique="DIVE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:25.80">
          <SWIMSTYLE distance="50" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:58.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="IMMERSION" technique="DIVE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:09:53.00">
          <SWIMSTYLE distance="800" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:04:40.00">
          <SWIMSTYLE distance="400" relaycount="1" stroke="IMMERSION" technique="DIVE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:08.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST name="Pflichtzeiten 2008 männlich" course="LCM" gender="M" timestandardlistid="23">
      <AGEGROUP agemax="15" agemin="15" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:04:45.00">
          <SWIMSTYLE distance="400" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:19:37.00">
          <SWIMSTYLE distance="1500" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:59.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:19:37.00">
          <SWIMSTYLE distance="1500" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:22.50">
          <SWIMSTYLE distance="50" relaycount="1" stroke="APNEA" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:10:04.00">
          <SWIMSTYLE distance="800" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:04:45.00">
          <SWIMSTYLE distance="400" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:04:50.00">
          <SWIMSTYLE distance="400" relaycount="1" stroke="IMMERSION" technique="DIVE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:26.30">
          <SWIMSTYLE distance="50" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:00.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="IMMERSION" technique="DIVE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:10:04.00">
          <SWIMSTYLE distance="800" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:04:50.00">
          <SWIMSTYLE distance="400" relaycount="1" stroke="IMMERSION" technique="DIVE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:10.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST name="Pflichtzeiten 2009 männlich" course="LCM" gender="M" timestandardlistid="24">
      <AGEGROUP agemax="14" agemin="14" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:04:55.00">
          <SWIMSTYLE distance="400" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:20:26.00">
          <SWIMSTYLE distance="1500" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:01.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:20:26.00">
          <SWIMSTYLE distance="1500" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:24.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="APNEA" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:10:24.00">
          <SWIMSTYLE distance="800" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:04:55.00">
          <SWIMSTYLE distance="400" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:05:04.00">
          <SWIMSTYLE distance="400" relaycount="1" stroke="IMMERSION" technique="DIVE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:27.10">
          <SWIMSTYLE distance="50" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:03.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="IMMERSION" technique="DIVE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:10:24.00">
          <SWIMSTYLE distance="800" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:05:04.00">
          <SWIMSTYLE distance="400" relaycount="1" stroke="IMMERSION" technique="DIVE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:15.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST name="Pflichtzeiten 2011 männlich" course="LCM" gender="M" timestandardlistid="25">
      <AGEGROUP agemax="12" agemin="12" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:21:26.00">
          <SWIMSTYLE distance="1500" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:21:26.00">
          <SWIMSTYLE distance="1500" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:11:10.00">
          <SWIMSTYLE distance="800" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:05:15.00">
          <SWIMSTYLE distance="400" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:05:15.00">
          <SWIMSTYLE distance="400" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:07.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:28.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="IMMERSION" technique="DIVE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:05:50.00">
          <SWIMSTYLE distance="400" relaycount="1" stroke="IMMERSION" technique="DIVE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:30.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:09.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="IMMERSION" technique="DIVE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:11:10.00">
          <SWIMSTYLE distance="800" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:05:50.00">
          <SWIMSTYLE distance="400" relaycount="1" stroke="IMMERSION" technique="DIVE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:30.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST name="Pflichtzeiten 2010 männlich" course="LCM" gender="M" timestandardlistid="26">
      <AGEGROUP agemax="13" agemin="13" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:20:56.00">
          <SWIMSTYLE distance="1500" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:20:56.00">
          <SWIMSTYLE distance="1500" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:10:40.00">
          <SWIMSTYLE distance="800" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:05:00.00">
          <SWIMSTYLE distance="400" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:05:00.00">
          <SWIMSTYLE distance="400" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:03.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:27.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="IMMERSION" technique="DIVE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:05:20.00">
          <SWIMSTYLE distance="400" relaycount="1" stroke="IMMERSION" technique="DIVE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:28.50">
          <SWIMSTYLE distance="50" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:05.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="IMMERSION" technique="DIVE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:10:40.00">
          <SWIMSTYLE distance="800" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:05:20.00">
          <SWIMSTYLE distance="400" relaycount="1" stroke="IMMERSION" technique="DIVE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:22.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST name="Pflichtzeiten 1959 bis 1968 männlich" course="LCM" gender="M" timestandardlistid="27">
      <AGEGROUP agemax="64" agemin="55" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:17:10.00">
          <SWIMSTYLE distance="1500" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:17:10.00">
          <SWIMSTYLE distance="1500" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST name="Pflichtzeiten 1959 bis 1968 weiblich" course="LCM" gender="F" timestandardlistid="28">
      <AGEGROUP agemax="64" agemin="55" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:17:50.00">
          <SWIMSTYLE distance="1500" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:17:50.00">
          <SWIMSTYLE distance="1500" relaycount="1" stroke="SURFACE" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
  </TIMESTANDARDLISTS>
</LENEX>
